# Spheral++ Visit dump file 1.1
# time  = 0
# cycle = 0
!Header
!Time 0
!Cycle 0
!NodeList "Earth"
!Field "position" Vector 3
!Field "gravitational_potential" Scalar 1
!Field "mass" Scalar 1
!Field "position" Vector 3
!Field "velocity" Vector 3
!Field "H" SymTensor 3 3
!Field "H_trace" Scalar 1
!Field "H_determinant" Scalar 1
!Field "H_eigen_min" Scalar 1
!Field "H_eigen_max" Scalar 1
!Field "work" Scalar 1
!Field "H_inverse" SymTensor 3 3
!Field "H_inverse_trace" Scalar 1
!Field "H_inverse_determinant" Scalar 1
!Field "H_inverse_eigen_min" Scalar 1
!Field "H_inverse_eigen_max" Scalar 1
!Field "hmin" Scalar 1
!Field "hmax" Scalar 1
!Field "hmin_hmax_ratio" Scalar 1
!Field "Domains" Scalar 1
!NodeList "fragments"
!Field "position" Vector 3
!Field "gravitational_potential" Scalar 1
!Field "mass" Scalar 1
!Field "position" Vector 3
!Field "velocity" Vector 3
!Field "H" SymTensor 3 3
!Field "H_trace" Scalar 1
!Field "H_determinant" Scalar 1
!Field "H_eigen_min" Scalar 1
!Field "H_eigen_max" Scalar 1
!Field "work" Scalar 1
!Field "H_inverse" SymTensor 3 3
!Field "H_inverse_trace" Scalar 1
!Field "H_inverse_determinant" Scalar 1
!Field "H_inverse_eigen_min" Scalar 1
!Field "H_inverse_eigen_max" Scalar 1
!Field "hmin" Scalar 1
!Field "hmax" Scalar 1
!Field "hmin_hmax_ratio" Scalar 1
!Field "Domains" Scalar 1
!EndHeader
!ASCIIData
!NodeList "Earth" 1
!Field "position" Vector 3
   -0.186807701696555666925903      0.98239649968169706628629                              0 
!Field "gravitational_potential" Scalar 1
                             0
!Field "mass" Scalar 1
3.002735152746214529484187e-06
!Field "position" Vector 3
   -0.186807701696555666925903      0.98239649968169706628629                              0 
!Field "velocity" Vector 3
    -6.17257925262469431260115    -1.173747406567785533937354                              0 
!Field "H" SymTensor 3 3
1.201671814746419312130462e-08                              0                              0                              0 1.201671814746419312130462e-08                              0                              0                              0 1.201671814746419312130462e-08 
!Field "H_trace" Scalar 1
3.605015444239258101827509e-08
!Field "H_determinant" Scalar 1
1.735232306249560992915282e-24
!Field "H_eigen_min" Scalar 1
1.201671814746419312130462e-08
!Field "H_eigen_max" Scalar 1
1.201671814746419312130462e-08
!Field "work" Scalar 1
0.0003999999999999999649585858
!Field "H_inverse" SymTensor 3 3
    83217396.60766059160232544                              0                              0                              0     83217396.60766059160232544                              0                              0                              0     83217396.60766059160232544 
!Field "H_inverse_trace" Scalar 1
    249652189.8229817748069763
!Field "H_inverse_determinant" Scalar 1
      576291714024935098679296
!Field "H_inverse_eigen_min" Scalar 1
    83217396.60766057670116425
!Field "H_inverse_eigen_max" Scalar 1
    83217396.60766057670116425
!Field "hmin" Scalar 1
    83217396.60766057670116425
!Field "hmax" Scalar 1
    83217396.60766057670116425
!Field "hmin_hmax_ratio" Scalar 1
                             1
!Field "Domains" Scalar 1
                             0
!NodeList "fragments" 100
!Field "position" Vector 3
  -0.1099958325213291343569466    0.7159336745622498776597809 -9.122899804995146994977612e-10 
  -0.1099958331352110796341748    0.7159336877092649098486277 -9.538393228485688617717299e-09 
  -0.1099958265342588364932297    0.7159336826645700257998328 9.325333913342428343804632e-10 
  -0.1099958305512364203915254    0.7159336768089165081718761 -4.621939848374083675230241e-09 
  -0.1099958309796880834285915    0.7159336758792127497486035 1.337943081372146478928642e-12 
  -0.1099958316281972048322757    0.7159336747698260561278971 7.560959482996491419114138e-10 
    -0.10999583178054934962109    0.7159336774073183917721508 5.166974015696412241985757e-09 
  -0.1099958310007940892605305    0.7159336759222961754645098 8.400549767855012441314019e-13 
  -0.1099958319441468601596057     0.715933676895159298858573  5.36745580805813947664671e-09 
  -0.1099958304172500428430581    0.7159336755049872103029429 -2.845204521125208339446122e-09 
  -0.1099958295233919164379799    0.7159336744400762730933252 -1.187906498672522982233374e-09 
  -0.1099958311142214956168672    0.7159336757870649048385303 -1.809746951606384688113895e-09 
  -0.1099958235931268318852361    0.7159336718917602704337355 7.405756417123649871579361e-09 
  -0.1099958308857647282241743    0.7159336758958492197280066 1.534439324506648843721797e-08 
  -0.1099958280457383336115029    0.7159336717868169941425549 -1.999044089618114261646652e-09 
  -0.1099958285785337247508764    0.7159336765482107178826254 4.521073201362273481612602e-10 
  -0.1099958294377303136268864    0.7159336761404488935767176 -7.265054344742333932976826e-10 
  -0.1099958301089067197464644    0.7159336771811330990544775 -9.889447015482376212343606e-10 
  -0.1099958314617641708110796    0.7159336715591969602101585   9.7242650922702875714774e-10 
  -0.1099958309492572311460989    0.7159336762707945167605317 -3.597396461795856625339801e-09 
  -0.1099958299863762894998942    0.7159336749147016121241904 -2.111596965830699906310307e-09 
  -0.1099958307655026779059426    0.7159336763550124826949173 8.961518935431247508662997e-10 
  -0.1099958351789761673567014    0.7159336763067569719964922 -1.863416206424479991117808e-09 
  -0.1099958295335490970900949    0.7159336859897665883423201 1.742003455891271359777486e-09 
  -0.1099958318026763720576255    0.7159336768556151531228693  -4.0770356372710929346248e-09 
  -0.1099958302913075641749074    0.7159336759382817216845751 7.989286235246487522274549e-10 
  -0.1099958302715921543146749    0.7159336757751525448512098  4.46615416718414080799201e-09 
  -0.1099958310682836865046497    0.7159336741689210636963026 -3.234496750253793017718404e-10 
  -0.1099958290748948436243992    0.7159336757346533852697235  -4.5482046671905180552769e-10 
  -0.1099958308925318289928086     0.715933675722448925604624 -1.990623560279041351167489e-10 
  -0.1099958297666315115703739    0.7159336753401355224468716 6.604192131845606517237195e-09 
  -0.1099958316739478580981171     0.715933675800253355170355 -4.122801568327054544098387e-09 
  -0.1099958308579942756200154    0.7159336761724892639335849 2.194155212619120340328058e-09 
  -0.1099958347252651402747858    0.7159336728313563380510232 -1.227265260178359600400771e-09 
  -0.1099958307173143912116586    0.7159336761496677414839951  -1.0023052818095029715283e-09 
  -0.1099958351569774450684491    0.7159336757884688928754713 -2.379518077207225043150225e-09 
  -0.1099958309875381234910208    0.7159336760497707619066432 4.051828198574202635388604e-11 
  -0.1099958305449326434466428    0.7159336771735036464292534 -2.189233992996437871301592e-09 
  -0.1099958381814055558001186    0.7159336822464633653950727 4.371996352786077348116164e-09 
  -0.1099958272376623524824168     0.715933679173659021088838 8.461002530228396915112004e-09 
    -0.10999583142596643103861    0.7159336770212707534710717 -1.679301275567199994522661e-09 
  -0.1099958312345346994609585    0.7159336698716022295840844 -1.592191061464689689051473e-08 
  -0.1099958316115887679842444    0.7159336752132318126840005 -4.908310688715580986523078e-10 
   -0.109995830210098885504344    0.7159336761653684044759416 8.079910030227324945916492e-09 
  -0.1099958233507539462348035     0.715933671264713966664317  3.06498034507972375434311e-09 
  -0.1099958300164498581352746    0.7159336743078057452294161 2.270254410036008094874274e-09 
  -0.1099958282504941986523761    0.7159336735750940761136007 5.077667640176801723916094e-10 
  -0.1099958309123191813050369    0.7159336758672152356552942 2.179496113256682668826123e-10 
  -0.1099958314929177366492397    0.7159336754272750402705583 5.516965913039183584502981e-09 
  -0.1099958310542294426248588    0.7159336753633637195903816 1.893580465287307013318677e-09 
  -0.1099958392777546645202591    0.7159336745479690788940275 1.226789279750542084293544e-10 
  -0.1099958309479215079473846    0.7159336783911638413258061 2.394287470002324491924126e-09 
  -0.1099958317169908994515026    0.7159336774239364320493451 -1.051086361067444997096384e-08 
  -0.1099958318814173025002034    0.7159336778838064629937321 -2.230048122572747255444343e-09 
  -0.1099958290221636353356516     0.715933678102552817357207 -5.395861021512033232138981e-09 
  -0.1099958301396516124892599    0.7159336776307195782109716 5.090286364558539958466454e-09 
  -0.1099958307152672093431889    0.7159336761345087563057632 2.204048544545941728334763e-10 
   -0.109995830501163474601789    0.7159336755012712938395225 1.591804197473800251273194e-09 
  -0.1099958309391784461173103    0.7159336758833410030433697 -5.285713289118255984055362e-11 
  -0.1099958378016106796959406    0.7159336773242274132300622 1.364968808958334562172393e-08 
  -0.1099958303176714197180175    0.7159336758104780651379428 3.213834392661391653672842e-10 
  -0.1099958325564137778806995    0.7159336798698145987174257 -3.270590002713228482905036e-09 
  -0.1099958299011249140963997    0.7159336752729030806108312 -1.726249855486896897836403e-09 
  -0.1099958245751296859182844    0.7159336781754910283837035 3.876489355986368048917336e-09 
  -0.1099958244033803905770341    0.7159336736405229606461376 6.306079982713442456963276e-09 
  -0.1099958213317608901604672     0.715933677439911098083769 2.742600630834892142973838e-09 
  -0.1099958338396684331961239    0.7159336823628207335801221 -5.527733972000049103752591e-09 
  -0.1099958335041015533573017    0.7159336733608520075833326 1.741155392451429394198727e-08 
  -0.1099958293919679475081352    0.7159336744927400353333269 2.651282500745213569348082e-09 
  -0.1099958326066814706667429    0.7159336722688557363980522 -4.355027415950067564494493e-09 
  -0.1099958311010877515245809    0.7159336734157225601293817 1.481107196440043362330305e-08 
  -0.1099958330774078313352149    0.7159336761920680469728495 -1.019009563524234560957292e-08 
  -0.1099958300925990839491675     0.715933676088634896039764 -3.665554570668681549094665e-09 
  -0.1099958339209717861351123     0.715933685228091976071596 5.910129821705691261507148e-10 
  -0.1099958283997590768876762    0.7159336657410794169109636 -6.021463484917284960179939e-09 
  -0.1099958319005117507449754    0.7159336728885590250825999  4.56821173111788490458234e-09 
   -0.109995835310012585184225    0.7159336786396820473399316 7.474913487591703169771948e-09 
  -0.1099958322954815576055765    0.7159336758937897560173269 6.702361159213309259407913e-09 
  -0.1099958210875019437580136    0.7159336785728641627812863 4.778817743820603432777138e-09 
  -0.1099958325544869858214625    0.7159336754998661955795569 -8.709509821160652344810822e-09 
  -0.1099958320778357118152613    0.7159336774463729291539948 1.124603449656185322869757e-08 
  -0.1099958294696939953283277    0.7159336752634788414439981 -3.407181803222010729685437e-09 
  -0.1099958338105815613960914    0.7159336762994249481195652 -1.931470912598449621680741e-09 
   -0.109995829937492128891563     0.715933677028878667769618 1.085738614309962985032451e-09 
  -0.1099958306834903920545798    0.7159336758561797298128226 7.218022214829826306396637e-10 
  -0.1099958307125486756117283     0.715933683126640296734422 -2.478595674483252380733595e-09 
  -0.1099958310694191532252972    0.7159336759949653794521396 6.169959217288334759526967e-09 
  -0.1099958305563912552837991     0.715933671578907970811656 -1.531463689545657607799075e-10 
  -0.1099958313444093088717679    0.7159336768321589161701013 -7.325658561314216190365118e-09 
   -0.109995837942509028239968    0.7159336778783700339090501 -4.631443168528082290571898e-09 
  -0.1099958197141485127801275    0.7159336693412646779322017 -9.33317565381944576576636e-09 
   -0.109995831662565560216116    0.7159336755115038863905852 -1.088963771310952616815792e-08 
   -0.109995832718991687348975    0.7159336750629933243672554 -8.061937756213157773881696e-10 
    -0.10999583207544130769584    0.7159336754924766621499543 -5.462138995734873966589553e-10 
  -0.1099958302518213026921501     0.715933674879680626013112 -3.196044722735010753162971e-10 
  -0.1099958308172675341962687    0.7159336762738194304134254 4.789318181641549975542685e-10 
  -0.1099958292524905734133256    0.7159336733569888755468469 -1.236485168538024533104166e-08 
  -0.1099958356024782618609592    0.7159336803413559602304872 -5.846170723618728431633251e-09 
  -0.1099958302182307695593622    0.7159336765051226292300157 -2.922412125294453445103358e-09 
   -0.109995830932486951536653    0.7159336759443410969083743 -3.858452492371351636233694e-10 
!Field "gravitational_potential" Scalar 1
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
!Field "mass" Scalar 1
1.730003566208363479963318e-21
1.124269785489431254374978e-21
1.329113979043533905521146e-21
1.254037367764818378525713e-21
1.062918052617490386895235e-21
1.895603121463646382377901e-23
3.533437029315092547222878e-22
1.510884874685156423995826e-21
3.021769859054850761975975e-21
2.882343673796532324218186e-21
9.807816975401448174789604e-22
1.072145875126913938149897e-21
7.363698323362288425709683e-22
7.882395196774288442180405e-22
 8.00876624778447601815496e-22
6.826319872878034312134189e-22
1.421645097437905637388497e-22
1.657220317410581502961611e-22
1.438785399582395571021306e-21
3.891004040471064309100272e-23
2.305738007096525332715661e-21
1.292863089421015571991463e-21
8.069131158595730315682619e-23
2.789228629298556340370964e-22
5.163614042843619635187599e-22
9.584246727593269365114201e-22
6.657736465745111485126499e-22
9.534152335076600231787535e-22
1.460971926760905966563326e-22
4.038166503514281151566608e-22
1.543443256323561530304135e-22
1.911416402774293614116787e-22
7.935942934874135286293355e-22
6.206920840176931468169757e-22
2.369226934796584631342291e-22
5.883657164556437259896445e-23
1.918827006107497457988563e-22
1.484499886919274691798193e-21
1.115734332452909752712497e-21
 2.16750070134820384593364e-21
1.827749799850109740128436e-22
3.404367993375842023846044e-22
2.907169574305044979063179e-21
7.431520000840151056281697e-23
3.032902264710393510379616e-22
2.244193331726852873018759e-21
2.606351393924481646614516e-21
5.714947496310070190279399e-22
8.460915786904154815108693e-23
8.253355763243080850631942e-22
 2.22364087818746642412756e-22
3.280910001636689996245908e-21
1.450868852173969275246061e-22
 2.26370326216586145402534e-21
1.213367416512781610964214e-22
4.748093171417177610473424e-23
1.976224611534000932611867e-21
9.221051052447671450131824e-22
3.035285472383758672026508e-23
3.382499899106131348140972e-22
2.987277232564295663511155e-22
6.401455058035773193497448e-23
1.105848699343182884780805e-22
8.727849596098254246973935e-22
5.765096068015846361555932e-22
1.628780775013538302893861e-21
 2.92217396070347831852402e-21
 1.53511423301234768365532e-22
3.569269987296214527359568e-22
5.796209110957019992751636e-22
4.449022433866837624611413e-22
1.119969811746083140979446e-22
3.459910725636516388309869e-22
4.676456605730311511545029e-22
1.170575647706002154792793e-21
8.539297151952041622468664e-22
4.976759339867310610258307e-22
1.605046839532581097117795e-21
8.974546492733593085165357e-22
5.533066247094537929008333e-22
1.777481078657949035729717e-21
1.249379440475242357419131e-21
2.357809191116508301206947e-22
4.237639998516635478710503e-22
9.226794695730891063046088e-22
2.199193805178737132092592e-21
9.092359064002320044819532e-22
3.991209002159260272071407e-22
6.057095919306659666940979e-22
4.228182669331054402224854e-22
1.046846517673758294402904e-21
9.785346942544565774757123e-22
3.144724265016950973472716e-22
1.262689223590133749672884e-21
4.355054974984577963817195e-22
3.115115652362280241118265e-21
2.004520908154835607507435e-22
8.642971912829557341333532e-23
2.691318063360457761827114e-22
5.983014467865911127126781e-22
!Field "position" Vector 3
  -0.1099958325213291343569466    0.7159336745622498776597809 -9.122899804995146994977612e-10 
  -0.1099958331352110796341748    0.7159336877092649098486277 -9.538393228485688617717299e-09 
  -0.1099958265342588364932297    0.7159336826645700257998328 9.325333913342428343804632e-10 
  -0.1099958305512364203915254    0.7159336768089165081718761 -4.621939848374083675230241e-09 
  -0.1099958309796880834285915    0.7159336758792127497486035 1.337943081372146478928642e-12 
  -0.1099958316281972048322757    0.7159336747698260561278971 7.560959482996491419114138e-10 
    -0.10999583178054934962109    0.7159336774073183917721508 5.166974015696412241985757e-09 
  -0.1099958310007940892605305    0.7159336759222961754645098 8.400549767855012441314019e-13 
  -0.1099958319441468601596057     0.715933676895159298858573  5.36745580805813947664671e-09 
  -0.1099958304172500428430581    0.7159336755049872103029429 -2.845204521125208339446122e-09 
  -0.1099958295233919164379799    0.7159336744400762730933252 -1.187906498672522982233374e-09 
  -0.1099958311142214956168672    0.7159336757870649048385303 -1.809746951606384688113895e-09 
  -0.1099958235931268318852361    0.7159336718917602704337355 7.405756417123649871579361e-09 
  -0.1099958308857647282241743    0.7159336758958492197280066 1.534439324506648843721797e-08 
  -0.1099958280457383336115029    0.7159336717868169941425549 -1.999044089618114261646652e-09 
  -0.1099958285785337247508764    0.7159336765482107178826254 4.521073201362273481612602e-10 
  -0.1099958294377303136268864    0.7159336761404488935767176 -7.265054344742333932976826e-10 
  -0.1099958301089067197464644    0.7159336771811330990544775 -9.889447015482376212343606e-10 
  -0.1099958314617641708110796    0.7159336715591969602101585   9.7242650922702875714774e-10 
  -0.1099958309492572311460989    0.7159336762707945167605317 -3.597396461795856625339801e-09 
  -0.1099958299863762894998942    0.7159336749147016121241904 -2.111596965830699906310307e-09 
  -0.1099958307655026779059426    0.7159336763550124826949173 8.961518935431247508662997e-10 
  -0.1099958351789761673567014    0.7159336763067569719964922 -1.863416206424479991117808e-09 
  -0.1099958295335490970900949    0.7159336859897665883423201 1.742003455891271359777486e-09 
  -0.1099958318026763720576255    0.7159336768556151531228693  -4.0770356372710929346248e-09 
  -0.1099958302913075641749074    0.7159336759382817216845751 7.989286235246487522274549e-10 
  -0.1099958302715921543146749    0.7159336757751525448512098  4.46615416718414080799201e-09 
  -0.1099958310682836865046497    0.7159336741689210636963026 -3.234496750253793017718404e-10 
  -0.1099958290748948436243992    0.7159336757346533852697235  -4.5482046671905180552769e-10 
  -0.1099958308925318289928086     0.715933675722448925604624 -1.990623560279041351167489e-10 
  -0.1099958297666315115703739    0.7159336753401355224468716 6.604192131845606517237195e-09 
  -0.1099958316739478580981171     0.715933675800253355170355 -4.122801568327054544098387e-09 
  -0.1099958308579942756200154    0.7159336761724892639335849 2.194155212619120340328058e-09 
  -0.1099958347252651402747858    0.7159336728313563380510232 -1.227265260178359600400771e-09 
  -0.1099958307173143912116586    0.7159336761496677414839951  -1.0023052818095029715283e-09 
  -0.1099958351569774450684491    0.7159336757884688928754713 -2.379518077207225043150225e-09 
  -0.1099958309875381234910208    0.7159336760497707619066432 4.051828198574202635388604e-11 
  -0.1099958305449326434466428    0.7159336771735036464292534 -2.189233992996437871301592e-09 
  -0.1099958381814055558001186    0.7159336822464633653950727 4.371996352786077348116164e-09 
  -0.1099958272376623524824168     0.715933679173659021088838 8.461002530228396915112004e-09 
    -0.10999583142596643103861    0.7159336770212707534710717 -1.679301275567199994522661e-09 
  -0.1099958312345346994609585    0.7159336698716022295840844 -1.592191061464689689051473e-08 
  -0.1099958316115887679842444    0.7159336752132318126840005 -4.908310688715580986523078e-10 
   -0.109995830210098885504344    0.7159336761653684044759416 8.079910030227324945916492e-09 
  -0.1099958233507539462348035     0.715933671264713966664317  3.06498034507972375434311e-09 
  -0.1099958300164498581352746    0.7159336743078057452294161 2.270254410036008094874274e-09 
  -0.1099958282504941986523761    0.7159336735750940761136007 5.077667640176801723916094e-10 
  -0.1099958309123191813050369    0.7159336758672152356552942 2.179496113256682668826123e-10 
  -0.1099958314929177366492397    0.7159336754272750402705583 5.516965913039183584502981e-09 
  -0.1099958310542294426248588    0.7159336753633637195903816 1.893580465287307013318677e-09 
  -0.1099958392777546645202591    0.7159336745479690788940275 1.226789279750542084293544e-10 
  -0.1099958309479215079473846    0.7159336783911638413258061 2.394287470002324491924126e-09 
  -0.1099958317169908994515026    0.7159336774239364320493451 -1.051086361067444997096384e-08 
  -0.1099958318814173025002034    0.7159336778838064629937321 -2.230048122572747255444343e-09 
  -0.1099958290221636353356516     0.715933678102552817357207 -5.395861021512033232138981e-09 
  -0.1099958301396516124892599    0.7159336776307195782109716 5.090286364558539958466454e-09 
  -0.1099958307152672093431889    0.7159336761345087563057632 2.204048544545941728334763e-10 
   -0.109995830501163474601789    0.7159336755012712938395225 1.591804197473800251273194e-09 
  -0.1099958309391784461173103    0.7159336758833410030433697 -5.285713289118255984055362e-11 
  -0.1099958378016106796959406    0.7159336773242274132300622 1.364968808958334562172393e-08 
  -0.1099958303176714197180175    0.7159336758104780651379428 3.213834392661391653672842e-10 
  -0.1099958325564137778806995    0.7159336798698145987174257 -3.270590002713228482905036e-09 
  -0.1099958299011249140963997    0.7159336752729030806108312 -1.726249855486896897836403e-09 
  -0.1099958245751296859182844    0.7159336781754910283837035 3.876489355986368048917336e-09 
  -0.1099958244033803905770341    0.7159336736405229606461376 6.306079982713442456963276e-09 
  -0.1099958213317608901604672     0.715933677439911098083769 2.742600630834892142973838e-09 
  -0.1099958338396684331961239    0.7159336823628207335801221 -5.527733972000049103752591e-09 
  -0.1099958335041015533573017    0.7159336733608520075833326 1.741155392451429394198727e-08 
  -0.1099958293919679475081352    0.7159336744927400353333269 2.651282500745213569348082e-09 
  -0.1099958326066814706667429    0.7159336722688557363980522 -4.355027415950067564494493e-09 
  -0.1099958311010877515245809    0.7159336734157225601293817 1.481107196440043362330305e-08 
  -0.1099958330774078313352149    0.7159336761920680469728495 -1.019009563524234560957292e-08 
  -0.1099958300925990839491675     0.715933676088634896039764 -3.665554570668681549094665e-09 
  -0.1099958339209717861351123     0.715933685228091976071596 5.910129821705691261507148e-10 
  -0.1099958283997590768876762    0.7159336657410794169109636 -6.021463484917284960179939e-09 
  -0.1099958319005117507449754    0.7159336728885590250825999  4.56821173111788490458234e-09 
   -0.109995835310012585184225    0.7159336786396820473399316 7.474913487591703169771948e-09 
  -0.1099958322954815576055765    0.7159336758937897560173269 6.702361159213309259407913e-09 
  -0.1099958210875019437580136    0.7159336785728641627812863 4.778817743820603432777138e-09 
  -0.1099958325544869858214625    0.7159336754998661955795569 -8.709509821160652344810822e-09 
  -0.1099958320778357118152613    0.7159336774463729291539948 1.124603449656185322869757e-08 
  -0.1099958294696939953283277    0.7159336752634788414439981 -3.407181803222010729685437e-09 
  -0.1099958338105815613960914    0.7159336762994249481195652 -1.931470912598449621680741e-09 
   -0.109995829937492128891563     0.715933677028878667769618 1.085738614309962985032451e-09 
  -0.1099958306834903920545798    0.7159336758561797298128226 7.218022214829826306396637e-10 
  -0.1099958307125486756117283     0.715933683126640296734422 -2.478595674483252380733595e-09 
  -0.1099958310694191532252972    0.7159336759949653794521396 6.169959217288334759526967e-09 
  -0.1099958305563912552837991     0.715933671578907970811656 -1.531463689545657607799075e-10 
  -0.1099958313444093088717679    0.7159336768321589161701013 -7.325658561314216190365118e-09 
   -0.109995837942509028239968    0.7159336778783700339090501 -4.631443168528082290571898e-09 
  -0.1099958197141485127801275    0.7159336693412646779322017 -9.33317565381944576576636e-09 
   -0.109995831662565560216116    0.7159336755115038863905852 -1.088963771310952616815792e-08 
   -0.109995832718991687348975    0.7159336750629933243672554 -8.061937756213157773881696e-10 
    -0.10999583207544130769584    0.7159336754924766621499543 -5.462138995734873966589553e-10 
  -0.1099958302518213026921501     0.715933674879680626013112 -3.196044722735010753162971e-10 
  -0.1099958308172675341962687    0.7159336762738194304134254 4.789318181641549975542685e-10 
  -0.1099958292524905734133256    0.7159336733569888755468469 -1.236485168538024533104166e-08 
  -0.1099958356024782618609592    0.7159336803413559602304872 -5.846170723618728431633251e-09 
  -0.1099958302182307695593622    0.7159336765051226292300157 -2.922412125294453445103358e-09 
   -0.109995830932486951536653    0.7159336759443410969083743 -3.858452492371351636233694e-10 
!Field "velocity" Vector 3
   -7.714378785873477362144968      4.23114101424258048922411 -8.540208487360047412135892e-06 
   -7.714366973261780557891143     4.231169597589506281565264 -1.310449826815465522000369e-05 
   -7.714352546250269782035502     4.231170924686009193749214 2.416120930159759252114698e-06 
   -7.714362233353718067974114     4.231157490028300216522439 -2.061209677867337122358221e-05 
   -7.714385037322768035039644     4.231153225300270825925963 6.583127853071149968285721e-07 
   -7.714373609630210459897626     4.231137846123004031539949 1.056084382183707289783962e-05 
    -7.71436721641701694807125     4.231159254672091307725168 1.998556131294559621625929e-05 
   -7.714381478426829197303505     4.231165083935596094022458 2.301895756211781949790505e-07 
   -7.714367778347035020658495     4.231157202223657876061225 2.038345789877549096998609e-05 
   -7.714360194701213480072965     4.231150636373024909175911 -2.057998406165663517913313e-05 
     -7.7143512168708223697422     4.231140375181649204705536 -1.070385819087819473393892e-05 
   -7.714366008123072937507914     4.231152274566029269919909 -2.096729907736289254672861e-05 
   -7.714350079010943161961222     4.231145811303988146789834 1.399119382945013399159682e-05 
   -7.714363882772817149202638     4.231153367524053798831574 2.109482377358110587054277e-05 
   -7.714352648189585437421556     4.231137341919009919877226 -7.816677486469657658578643e-06 
   -7.714343994868054998903517     4.231159004601417805702113  3.82614564154418855540388e-06 
   -7.714345198562448047141515     4.231156610113186999910795 -9.088874532405981905114171e-06 
   -7.714354421907854586493158     4.231168329810944150892738 -1.138466821488332293677535e-05 
     -7.7143664361537975793226     4.231132908003352177672696 4.600063288735828567201872e-06 
    -7.71436402539039889347805     4.231155626304531125470021 -2.097110814597448520831512e-05 
   -7.714355960444407855902682      4.23114523224717764549041 -1.775668268423057172896058e-05 
    -7.71436044015857191880059     4.231163095225562997825364  1.83736206952918476825818e-05 
   -7.714383185141323373557043     4.231155282198358236200875 -8.447980760678159913739695e-06 
   -7.714361094189905010409802     4.231173941834763141400799 3.548830578922066064423337e-06 
   -7.714368219728664932688389     4.231158155371340434669492 -2.009109569734170131459494e-05 
   -7.714350716942587560254196      4.23115455116027927573441 1.638137274911450415358985e-05 
   -7.714360845956377055188113     4.231152857837507497151819 2.085919676931753289706242e-05 
   -7.714365541290185035450122     4.231132676185963781279042 -3.908319526396067756580151e-06 
   -7.714343518785724107544866     4.231151755826306981589369 -4.991504947711142426553226e-06 
   -7.714360321622413252384831     4.231140476196469712988346 -1.631577333403580468075729e-05 
   -7.714360284316034821472385     4.231151654182998100850455 2.070456667281925805675601e-05 
   -7.714367664992381357080831     4.231152946131854442057829 -2.076195892037688018596717e-05 
   -7.714363202128241780997087     4.231156135692321740293664 2.089605724684469328531963e-05 
   -7.714379888820414699068806     4.231140523307671763575399 -5.162430297403541752654637e-06 
   -7.714359588604029482894475     4.231158717138665537049746 -1.992709718690877649435039e-05 
   -7.714382324995324502481253     4.231152948882997755220003 -1.03590222219562039289659e-05 
   -7.714369821153736594965267     4.231173057154663297296793 4.689570904468185895581922e-06 
    -7.71436074006399330471595     4.231163953891359241765713 -1.794785018047342518691424e-05 
   -7.714378384661443099901135     4.231166028501802678363219 8.709315971311383928923737e-06 
   -7.714355993830154467616467      4.23116043280415254912441 1.820471766192622455993004e-05 
   -7.714368892768572294471596      4.23116487632067617141729 -1.695947850016765189626149e-05 
   -7.714364321951458158821424     4.231145898850214415176652 -1.973362441784023402191993e-05 
   -7.714377283867230872260734     4.231140182588278619846278 -9.697207832663207866235461e-06 
   -7.714362064425232645703545     4.231154087982277545165744 2.099710291030481228808854e-05 
   -7.714346917015960869434821     4.231142981720506845988439 6.882986947010531349438849e-06 
   -7.714357282226933065771846     4.231141954018202255838332 1.645429564420771199016735e-05 
   -7.714348104028331043480193     4.231139749650422388072002  2.99573611491933006358403e-06 
   -7.714361598519653639982607     4.231152169480866476192205 2.093016264024953246693575e-05 
   -7.714366061525554485456269      4.23115163041331143745083 2.091916148964530604509662e-05 
    -7.71436521249385354082051     4.231147807823299800134009 2.031626141057306540998323e-05 
   -7.714384781991770800857466     4.231150019987517829633816 3.063548039354607445023683e-07 
   -7.714364020370372720947216     4.231168613930382349508363 1.455513192348664802081449e-05 
   -7.714365497933085791260055     4.231156403540337507251934 -2.081478836261393042098879e-05 
   -7.714370291364730292116292     4.231166794697196031904696 -1.496419949818579614626585e-05 
    -7.71435737689841705133631      4.23116098037759957861681 -1.853248329841529707046402e-05 
   -7.714360862737005497535847     4.231160133671699519197773 1.973223666391863629818691e-05 
   -7.714352366180682984975192     4.231166682775129750382348  1.15259023783361814406408e-05 
   -7.714358524855850163248761     4.231148633117808977033292 1.983256751224802009927334e-05 
   -7.714364884156709400997443     4.231154889789634054864109 -2.10176956756763355226459e-05 
   -7.714373388919278262676471     4.231155330889432519825277 1.876209882662779719359608e-05 
   -7.714345320844126163706278     4.231151269278830895359533  9.67118466046502244957625e-06 
   -7.714370270860049672023706     4.231168911143021738041625 -1.275838044782132339152909e-05 
   -7.714353561451753549249588       4.2311472593032810607383 -1.73198593390883302529492e-05 
   -7.714346737998850400686024     4.231159558132642217742614 1.048990599037002386197982e-05 
   -7.714349216187032176605953      4.23114829487281962627776 1.422392969292663288528693e-05 
   -7.714343911799403485929361     4.231156600908485998502329 5.722491713063592439609227e-06 
   -7.714370756200015222248112     4.231168539711640974587681 -1.29550622433258588690275e-05 
   -7.714366999051303075418673      4.23115035665668948183793 2.065885726638030708813241e-05 
   -7.714354275005240069162937     4.231144657771354289366172 1.660921510535741168687607e-05 
   -7.714369924996928418181596     4.231140432080719548935122 -1.557526679337750978495553e-05 
   -7.714364183737392188788817     4.231149883738009265243818 2.080777579772862562212422e-05 
   -7.714368287670886559226346     4.231153978031111151381083 -2.063508603694302694607499e-05 
    -7.71435922572482102310687     4.231154516272499499507376 -2.052506117205259606340456e-05 
   -7.714370356125423100479566     4.231173404613470800939012 1.268152860616575063716096e-06 
   -7.714359515789809940145005     4.231135613582692300838062 -1.053117378269492789553442e-05 
   -7.714367619370788631272262     4.231141965857436737508124 1.738016226904487017521257e-05 
    -7.71437410234223630567385     4.231159750977515621173097 1.734793509024343174246274e-05 
   -7.714368143922037290849403     4.231153389201901759975044 2.067440722014522732990181e-05 
   -7.714345523589751785209501     4.231158384706606767622361 8.941793580566677419256376e-06 
   -7.714367801617464159846804     4.231152441886186998942776 -2.072123208164315945572879e-05 
   -7.714366062135253443443617     4.231156241452724842133648 2.078843424469167949233082e-05 
   -7.714355722724398845002725     4.231149889527780594278283 -1.911333691574820093208101e-05 
   -7.714381333562658760172326     4.231155884984261206227529 -1.168164973940266358515445e-05 
   -7.714352682539901806535454     4.231166307988605268519677 1.224478289286281766483095e-05 
   -7.714356969915293404937984     4.231152703415615334847644 1.989527984152588289327827e-05 
    -7.71436333552487152331878     4.231173296313484044617326 -6.823514986798399618818031e-06 
   -7.714364406096967385906282     4.231153739751047027084496 2.108639082843139007819415e-05 
   -7.714362095260064222657093      4.23113234530503756758435 -7.478175044932797290041693e-07 
   -7.714365115061699640364168     4.231156061348396946186767 -2.088702914389509998150177e-05 
   -7.714381071902361775016743     4.231158229492880451516612 -1.131729999179845699874055e-05 
   -7.714349150961540502180469     4.231144721522468010732609 -1.230987416895537944565818e-05 
    -7.71436535492798647339896     4.231152634187320238368102 -2.103631015502801664173241e-05 
   -7.714381689708313061260014     4.231145219222291586902429 -8.023564834245797792598894e-06 
   -7.714382137977263020900409     4.231147164425479445526435 -8.723744324919771337290691e-06 
   -7.714352423801472902198384     4.231136518221187081678636  -5.3791180104981398536583e-06 
   -7.714359960850905473250805     4.231166511860681822554398 1.599041415407415151687769e-05 
   -7.714361162159681484240537     4.231149165464183070639592 -2.048755503810491593709789e-05 
   -7.714375253527727238633815     4.231164152052765636824461 -1.415987584083881013546566e-05 
   -7.714359021343573097340141     4.231157638805600917919492 -2.00558986766770914306722e-05 
   -7.714363718484526621921304     4.231156843053716976044143 -2.080157612070897315192583e-05 
!Field "H" SymTensor 3 3
1.201671814743165018164556e-08 7.193493479006149871751719e-20 6.297367362396827340179778e-20 7.193493479006149871751719e-20 1.201671814741524553573741e-08 -3.949373834634430633673541e-21 6.297367362396827340179778e-20 -3.949373834634430633673541e-21 1.201671814754567702908599e-08 
1.206246832727069008614682e-08 -1.261247774893291712398555e-19 7.762821215111084994673837e-20 -1.261247774893291712398555e-19  1.20624683279781561573675e-08 -3.281719656103199956681754e-19 7.762821215111084994673837e-20 -3.281719656103199956681754e-19 1.206246832782455864378375e-08 
1.206246832763782262049991e-08 1.976308191317819251079518e-19 1.015595812480356318653618e-19 1.976308191317819251079518e-19 1.206246832782142362926218e-08 1.463737452943210122068701e-20 1.015595812480356318653618e-19 1.463737452943210122068701e-20 1.206246832761390552026855e-08 
1.201671814732099326802067e-08 -3.14047391361882487041679e-20 -1.108690854520136818322021e-20 -3.14047391361882487041679e-20 1.201671814735184214178522e-08 -6.440562666187413343545955e-20 -1.108690854520136818322021e-20 -6.440562666187413343545955e-20 1.201671814771988953789579e-08 
1.201671814739731556877971e-08 -9.064245152356077261240896e-21 6.454283524598136690102884e-20 -9.064245152356077261240896e-21  1.20167181473901455672301e-08 -1.461731539957769029957138e-20 6.454283524598136690102884e-20 -1.461731539957769029957138e-20 1.201671814760529524455514e-08 
 1.20167181473909032646712e-08 5.013624410745156040163095e-20 5.213822798498302563173848e-21 5.013624410745156040163095e-20 1.201671814740540870389293e-08 -2.007401910543687561377935e-20 5.213822798498302563173848e-21 -2.007401910543687561377935e-20 1.201671814759635011341099e-08 
1.206246832756607462852828e-08 -8.669597282107027757559747e-20 -4.883612297967133915365182e-20 -8.669597282107027757559747e-20 1.206246832758197469426278e-08 1.016494337420742044965447e-19 -4.883612297967133915365182e-20 1.016494337420742044965447e-19 1.206246832792524637666616e-08 
1.201671814739997578162968e-08 -8.160963923448171040281318e-21 6.762739175019160710062432e-20 -8.160963923448171040281318e-21 1.201671814739026798996076e-08 -1.622173559520085660344384e-20 6.762739175019160710062432e-20 -1.622173559520085660344384e-20 1.201671814760250764589084e-08 
1.206246832759088177509875e-08 -6.983224167295170236799406e-20 -5.71663487359631734819037e-20 -6.983224167295170236799406e-20 1.206246832752546667789683e-08 6.031242679823204511481774e-20 -5.71663487359631734819037e-20 6.031242679823204511481774e-20 1.206246832795689761562489e-08 
1.201671814735332610380414e-08 -5.834683886765291310240455e-20 -5.960482548298121450319493e-22 -5.834683886765291310240455e-20 1.201671814736793080469937e-08 -3.100938557747911489875163e-21 -5.960482548298121450319493e-22 -3.100938557747911489875163e-21 1.201671814767144322377978e-08 
1.206246832761768904439037e-08 -1.349702333696649726810929e-19 -1.066184110792568108679566e-20 -1.349702333696649726810929e-19 1.206246832767135155944913e-08 3.050838554491047408998537e-20 -1.066184110792568108679566e-20 3.050838554491047408998537e-20 1.206246832778420877350342e-08 
1.201671814737190458036208e-08 -2.964780751512561792274103e-20 2.321747345420030561203716e-20 -2.964780751512561792274103e-20 1.201671814738068758410617e-08 -3.160119453166959277694986e-20 2.321747345420030561203716e-20 -3.160119453166959277694986e-20 1.201671814764022873618448e-08 
 1.20624683277609865049866e-08 -2.27516027482710261973381e-19 1.898331425936093869096281e-19 -2.27516027482710261973381e-19 1.206246832748688035668246e-08 -1.420486246664343687518862e-19 1.898331425936093869096281e-19 -1.420486246664343687518862e-19 1.206246832782547185118001e-08 
1.206246832745617706670571e-08 -2.682836239723862309294183e-20 -1.531879040841680004997718e-20 -2.682836239723862309294183e-20 1.206246832738681300925947e-08 -1.885692623164166451866543e-20 -1.531879040841680004997718e-20 -1.885692623164166451866543e-20 1.206246832823016831151036e-08 
1.206246832759840415558931e-08 -2.492121477693636248575831e-19 4.296169306447287486363379e-21 -2.492121477693636248575831e-19 1.206246832774579285149523e-08 8.342985017240464780136772e-20 4.296169306447287486363379e-21 8.342985017240464780136772e-20 1.206246832772920457149109e-08 
1.201671814751310596528611e-08  5.55695799610061226840238e-20 6.518875990680871238664405e-20  5.55695799610061226840238e-20 1.201671814734463078120498e-08 -2.071467048985919554796725e-20 6.518875990680871238664405e-20 -2.071467048985919554796725e-20 1.201671814753487570464728e-08 
1.201671814746651915318712e-08                              0                              0                              0 1.201671814734793950365519e-08                              0                              0                              0  1.20167181475781703379083e-08 
1.201671814736199826534614e-08 3.903465310637737597718178e-20 2.395122143162605458282036e-20 3.903465310637737597718178e-20 1.201671814744919137371536e-08 -3.921135956473401651422618e-20 2.395122143162605458282036e-20 -3.921135956473401651422618e-20 1.201671814758183805674436e-08 
1.206246832749329762387464e-08 5.214980851355876801918668e-20 1.880657161185249895895763e-20 5.214980851355876801918668e-20 1.206246832786083878545033e-08 -3.149844318995402137046193e-20 1.880657161185249895895763e-20 -3.149844318995402137046193e-20 1.206246832771899550837096e-08 
1.201671814734537193503383e-08 -4.845872182519402027699174e-20 2.990743882989069948419129e-20 -4.845872182519402027699174e-20 1.201671814736075749442731e-08 -5.471380991853173099013965e-20 2.990743882989069948419129e-20 -5.471380991853173099013965e-20 1.201671814768659220951808e-08 
1.201671814737065057455345e-08 -9.193285327914349578520836e-20 -1.488987141141391291844151e-20 -9.193285327914349578520836e-20 1.201671814739872177582105e-08 4.775137900388461248651732e-20 -1.488987141141391291844151e-20 4.775137900388461248651732e-20 1.201671814762328973160062e-08 
1.201671814737634157716781e-08 -3.012178200611850278044235e-20 4.775954741243357363480668e-20 -3.012178200611850278044235e-20 1.201671814737906465574434e-08 1.024690663315376857938829e-20 4.775954741243357363480668e-20 1.024690663315376857938829e-20 1.201671814763721118130989e-08 
1.206246832784378397558071e-08 -4.595939560436504715736777e-20 8.322039253166973582482137e-20 -4.595939560436504715736777e-20 1.206246832750154130585935e-08 1.228735440916894959637734e-20 8.322039253166973582482137e-20 1.228735440916894959637734e-20 1.206246832772788108251101e-08 
1.206246832742665995372737e-08   7.2545600877278771398491e-20 6.508381136659104700039474e-20   7.2545600877278771398491e-20 1.206246832800704130435785e-08 8.916965644291010683730042e-20 6.508381136659104700039474e-20 8.916965644291010683730042e-20 1.206246832763948856225359e-08 
1.201671814733275577633117e-08 -5.51282791042090824194799e-20 7.784886257950937007901032e-20 -5.51282791042090824194799e-20 1.201671814737855511248701e-08 -5.847867077777855188808719e-20 7.784886257950937007901032e-20 -5.847867077777855188808719e-20 1.201671814768153648161415e-08 
1.201671814739589943557102e-08 -4.40390958123231934101538e-21 6.303405780868464442206339e-20 -4.40390958123231934101538e-21 1.201671814736979030671639e-08 -1.805704257930288675706477e-20 6.303405780868464442206339e-20 -1.805704257930288675706477e-20 1.201671814762698226585506e-08 
1.206246832757576091350128e-08 -4.204476335545784368603883e-20 3.413786989585989576725288e-20 -4.204476335545784368603883e-20 1.206246832753404288648778e-08 -1.969948723370935005186648e-20 3.413786989585989576725288e-20 -1.969948723370935005186648e-20 1.206246832796360274167024e-08 
1.201671814734109210254448e-08 4.277428495694132953104574e-21 3.505136486662827120883851e-20 4.277428495694132953104574e-21 1.201671814749986942112403e-08 6.423458122083465268156504e-21 3.505136486662827120883851e-20 6.423458122083465268156504e-21 1.201671814755172371936376e-08 
1.201671814752495450038032e-08 -5.933904201241026979841281e-20 1.156222720468965171089319e-20 -5.933904201241026979841281e-20 1.201671814734220879637143e-08 -2.565562708379156810689289e-20 1.156222720468965171089319e-20 -2.565562708379156810689289e-20 1.201671814752558315764586e-08 
1.201671814738804783719666e-08 -1.383294138372428180687457e-20 4.178916454617895813450357e-20 -1.383294138372428180687457e-20 1.201671814739057900987108e-08  -6.4758936181010845381089e-21 4.178916454617895813450357e-20  -6.4758936181010845381089e-21 1.201671814761411298988496e-08 
 1.20624683275932905250425e-08 -6.128912030650403254192216e-20 5.660845418688736973837519e-20 -6.128912030650403254192216e-20 1.206246832748188253142141e-08 -3.714423521396400035472253e-20 5.660845418688736973837519e-20 -3.714423521396400035472253e-20 1.206246832799812098863208e-08 
1.201671814734316170843709e-08 -2.442912503052856632197731e-20 6.618065285883636169727423e-20 -2.442912503052856632197731e-20 1.201671814735186199411992e-08 -1.036126435283922465543927e-20 6.618065285883636169727423e-20 -1.036126435283922465543927e-20 1.201671814769780712426307e-08 
1.201671814734244206130417e-08 -3.437679907709127713998087e-20 1.678576937538545234924678e-20 -3.437679907709127713998087e-20 1.201671814735855057655302e-08 2.329650797679033317815964e-20 1.678576937538545234924678e-20 2.329650797679033317815964e-20  1.20167181476916347025322e-08 
1.206246832772079379902265e-08 1.766824701188764992418334e-19 7.546513484928468257694964e-20 1.766824701188764992418334e-19 1.206246832765089207417825e-08 1.359781529460608369029237e-20 7.546513484928468257694964e-20 1.359781529460608369029237e-20 1.206246832770165614837063e-08 
1.201671814738239819361293e-08 -1.104120681635781340418356e-20 3.485263472446240630995065e-20 -1.104120681635781340418356e-20 1.201671814739052607031187e-08 -3.747329800139525167663231e-20 3.485263472446240630995065e-20 -3.747329800139525167663231e-20 1.201671814762000913329123e-08 
1.206246832783284699352154e-08   4.5810813286835209561269e-21 1.030021842363281121303376e-19   4.5810813286835209561269e-21 1.206246832750232712744127e-08 1.050757192368454142543215e-20 1.030021842363281121303376e-19 1.050757192368454142543215e-20 1.206246832773811330668829e-08 
1.201671814739433275549084e-08 -2.161836530907337828276427e-20 3.388076374378508838989602e-20 -2.161836530907337828276427e-20 1.201671814738300203546009e-08 -2.598784268951461090049703e-20 3.388076374378508838989602e-20 -2.598784268951461090049703e-20 1.201671814761559529754265e-08 
1.201671814734149742104463e-08                              0                              0                              0 1.201671814743283635864396e-08 -6.805008104320620424248361e-20                              0 -6.805008104320620424248361e-20 1.201671814761831672175795e-08 
1.206246832772484698402416e-08 -3.275436702362976865848809e-19 -1.345618129422169152666251e-19 -3.275436702362976865848809e-19 1.206246832761224950468222e-08 8.515214360531662054890935e-20 -1.345618129422169152666251e-19 8.515214360531662054890935e-20 1.206246832773622402616922e-08 
1.206246832760480818789169e-08 9.707460796677311581220904e-20 1.403769960460412689494305e-19 9.707460796677311581220904e-20 1.206246832753800342726068e-08 1.288319328390620925627909e-19 1.403769960460412689494305e-19 1.288319328390620925627909e-19 1.206246832793048242994362e-08 
 1.20167181473863372276899e-08 -7.676732392859628639411596e-20 5.202976392716200987787097e-20 -7.676732392859628639411596e-20 1.201671814742536360899016e-08 -7.19665615237945808850236e-20 5.202976392716200987787097e-20 -7.19665615237945808850236e-20 1.201671814758099102379711e-08 
1.206246832733553442872608e-08 -8.096195681485268973338887e-20  6.10186322461991924922392e-20 -8.096195681485268973338887e-20 1.206246832754029802627991e-08 3.276977326253856879893257e-19  6.10186322461991924922392e-20 3.276977326253856879893257e-19 1.206246832819746324445124e-08 
 1.20167181474171033833932e-08 2.386498785276740144771501e-20  5.17585520838211859289725e-20 2.386498785276740144771501e-20 1.201671814739768945441658e-08 -6.427193359537025033750846e-21  5.17585520838211859289725e-20 -6.427193359537025033750846e-21 1.201671814757789736830616e-08 
1.206246832756995906868483e-08 -4.320984724823878316609521e-20  3.04281167137501525528793e-20 -4.320984724823878316609521e-20 1.206246832744570330578957e-08 -3.483722848555360616950617e-21  3.04281167137501525528793e-20 -3.483722848555360616950617e-21 1.206246832805778221749308e-08 
 1.20624683277948893295727e-08 -2.82611219362417223285866e-19 1.496113302118535625263168e-19 -2.82611219362417223285866e-19 1.206246832758306657267135e-08 -1.353515636320519184392086e-20 1.496113302118535625263168e-19 -1.353515636320519184392086e-20 1.206246832769534310593562e-08 
1.201671814734323780905344e-08 -7.982954655626759484648991e-20 6.004772900221507625885889e-20 -7.982954655626759484648991e-20 1.201671814742052791112917e-08 -7.350208015933149421179075e-20 6.004772900221507625885889e-20 -7.350208015933149421179075e-20 1.201671814762894764699048e-08 
1.206246832764751386855658e-08 -1.596301417910958337243593e-19 8.117019953406291445053775e-20 -1.596301417910958337243593e-19 1.206246832762472669704197e-08 4.738504139010019035500865e-21 8.117019953406291445053775e-20 4.738504139010019035500865e-21 1.206246832780101873791172e-08 
 1.20167181473811309529145e-08 -1.11818275204918281089117e-20 4.183197114287857731667816e-20 -1.11818275204918281089117e-20 1.201671814738943584626453e-08 -4.702521782363962331643958e-21 4.183197114287857731667816e-20 -4.702521782363962331643958e-21  1.20167181476222276316941e-08 
1.201671814732753792102719e-08 -1.604482234169107780948071e-20 -5.369911780087058885422083e-20 -1.604482234169107780948071e-20 1.201671814732343841391137e-08 -4.012859946647875507719921e-20 -5.369911780087058885422083e-20 -4.012859946647875507719921e-20  1.20167181477418528375203e-08 
1.201671814735651736660737e-08                              0                              0                              0 1.201671814736330355635275e-08 -2.851519046138738477892335e-20                              0 -2.851519046138738477892335e-20 1.201671814767321835337432e-08 
1.206246832799899283699771e-08 1.099984778573016202043999e-19 -1.499393460988220514225756e-20 1.099984778573016202043999e-19 1.206246832740692342431186e-08 -5.062203177156746818581403e-21 -1.499393460988220514225756e-20 -5.062203177156746818581403e-21 1.206246832766735131400683e-08 
1.206246832751186121118156e-08 -4.418467960013252628093117e-20 2.131272207273503455689928e-20 -4.418467960013252628093117e-20 1.206246832771309936496468e-08 8.497497185786541893379783e-20 2.131272207273503455689928e-20 8.497497185786541893379783e-20   1.2062468327848283838113e-08 
1.206246832740697470950983e-08 -7.356117187434075112631437e-20 4.115089130601772815488092e-20 -7.356117187434075112631437e-20 1.206246832756439048880113e-08 -7.856947906471083973545494e-20 4.115089130601772815488092e-20 -7.856947906471083973545494e-20 1.206246832810197186017689e-08 
 1.20167181473597350991902e-08 -1.119489697417016594617467e-19 5.254651916546037163563204e-20 -1.119489697417016594617467e-19 1.201671814747921637558981e-08 -7.950177623854345763032211e-20 5.254651916546037163563204e-20 -7.950177623854345763032211e-20 1.201671814755377347292166e-08 
1.201671814737001033675933e-08 6.167127774950353132771275e-20 -1.069188973614637693119111e-19 6.167127774950353132771275e-20 1.201671814738017307776516e-08 -1.152851313237958026261347e-19 -1.069188973614637693119111e-19 -1.152851313237958026261347e-19 1.201671814764243399969755e-08 
1.201671814733991254299098e-08  8.40534409566930615397614e-21 3.742082373128641898350766e-20  8.40534409566930615397614e-21 1.201671814735366855657774e-08 8.175935892535380841196491e-20 3.742082373128641898350766e-20 8.175935892535380841196491e-20 1.201671814769929604936567e-08 
1.201671814740074009651568e-08 -4.803851407401708221815706e-21 5.288460339144727941562089e-20 -4.803851407401708221815706e-21 1.201671814737569968501247e-08 -3.152385314439588468934939e-21 5.288460339144727941562089e-20 -3.152385314439588468934939e-21 1.201671814761640593454295e-08 
1.201671814736388589150399e-08 -3.213844833952278425177884e-20 5.120392748310438087297122e-20 -3.213844833952278425177884e-20 1.201671814736690510073981e-08 -3.216279846880481400395787e-20 5.120392748310438087297122e-20 -3.216279846880481400395787e-20 1.201671814766186943537009e-08 
1.201671814740312403104106e-08 -6.125272435955169932422781e-21  5.30090746865909033691029e-20 -6.125272435955169932422781e-21 1.201671814737798601222557e-08 -1.058142364274904142752926e-20  5.30090746865909033691029e-20 -1.058142364274904142752926e-20 1.201671814761175387077796e-08 
1.206246832769396502303511e-08 -1.431849640329290905202408e-19 -2.882790609196305689140849e-19 -1.431849640329290905202408e-19 1.206246832728446264334583e-08 1.947389957102965403566014e-21 -2.882790609196305689140849e-19 1.947389957102965403566014e-21 1.206246832809478862373748e-08 
1.201671814740201230029778e-08 -2.054964795765486652683041e-20 6.654688707504421470032355e-20 -2.054964795765486652683041e-20 1.201671814738594018099588e-08 2.272678732989443536709195e-21 6.654688707504421470032355e-20 2.272678732989443536709195e-21 1.201671814760473607046106e-08 
1.206246832751301264659423e-08 -1.289272654046588290023198e-19 7.409718491127511305963105e-20 -1.289272654046588290023198e-19 1.206246832779051023540985e-08 -1.031945037287466910647452e-19 7.409718491127511305963105e-20 -1.031945037287466910647452e-19 1.206246832776976950873069e-08 
1.201671814739810139036163e-08 -7.570522402207819885958107e-20 -1.377715839116523700305043e-20 -7.570522402207819885958107e-20 1.201671814737216596943565e-08 2.285830904729036676739651e-20 -1.377715839116523700305043e-20 2.285830904729036676739651e-20 1.201671814762249067512889e-08 
1.206246832785491782662568e-08 1.214325954646221217541474e-19 1.363522453780879436688843e-19 1.214325954646221217541474e-19 1.206246832751141784237323e-08 3.773577274951598427071495e-20 1.363522453780879436688843e-19 3.773577274951598427071495e-20 1.206246832770708245318897e-08 
1.206246832778996098748311e-08 -1.518761507290237523001147e-19 1.867516944790447561343421e-19 -1.518761507290237523001147e-19 1.206246832746663759273206e-08 -7.350519501132563920662894e-20 1.867516944790447561343421e-19 -7.350519501132563920662894e-20 1.206246832781653499184199e-08 
1.206246832799892666254871e-08 8.797810277052747047164816e-20 1.112471069919504154796183e-19 8.797810277052747047164816e-20 1.206246832743004643115516e-08 -1.502883775432282156781991e-20 1.112471069919504154796183e-19 -1.502883775432282156781991e-20 1.206246832764412904549001e-08 
1.206246832746454978886598e-08 -1.687721419210318955870381e-19 1.131874659138466801479479e-19 -1.687721419210318955870381e-19 1.206246832782606245813738e-08 -1.611749015850386129071817e-19 1.131874659138466801479479e-19 -1.611749015850386129071817e-19 1.206246832778266360011917e-08 
 1.20624683274379956368418e-08 -2.711001739581292901623555e-20 -1.655738480825956140821478e-19 -2.711001739581292901623555e-20 1.206246832736253360391981e-08 -1.87955287506749160394981e-19 -1.655738480825956140821478e-19 -1.87955287506749160394981e-19 1.206246832827270855605273e-08 
 1.20624683275971120994725e-08 -9.583714577039378641060141e-20 8.549893907712947740159919e-20 -9.583714577039378641060141e-20 1.206246832760258968948882e-08 -4.772439223640006995862464e-20 8.549893907712947740159919e-20 -4.772439223640006995862464e-20 1.206246832787337057173051e-08 
1.206246832751642890252408e-08 7.126533208419982281470878e-20 9.420346406060155675273038e-20 7.126533208419982281470878e-20 1.206246832773766166607383e-08 1.441412882186169596408516e-19 9.420346406060155675273038e-20 1.441412882186169596408516e-19 1.206246832781915715438378e-08 
1.206246832743594753764512e-08 -6.321893267559024610739715e-20 -4.270919618249106316587929e-20 -6.321893267559024610739715e-20 1.206246832743561997412255e-08 -1.507681422985089717296245e-19 -4.270919618249106316587929e-20 -1.507681422985089717296245e-19  1.20624683282019349828427e-08 
 1.20624683274645580606721e-08 -6.975365951475916473888128e-20 1.326493713659943152823224e-19 -6.975365951475916473888128e-20 1.206246832752093538250127e-08 1.720060045258079572819479e-20 1.326493713659943152823224e-19 1.720060045258079572819479e-20 1.206246832808788166562266e-08 
1.201671814736216701019111e-08 -4.914859045606324535783449e-20 -3.252081257767542129448815e-20 -4.914859045606324535783449e-20  1.20167181473394195433459e-08 -7.715423766011796508903706e-21 -3.252081257767542129448815e-20 -7.715423766011796508903706e-21 1.201671814769115659213815e-08 
1.206246832745723420352856e-08 -1.969289563820306811258234e-19 7.559913810851827306027881e-21 -1.969289563820306811258234e-19 1.206246832796472108985841e-08 2.546317834440227776191109e-20 7.559913810851827306027881e-21 2.546317834440227776191109e-20 1.206246832765136853021108e-08 
1.206246832739452398692969e-08 -1.856863310865162054828087e-19 -6.480960099352971832617487e-21 -1.856863310865162054828087e-19 1.206246832798817496894674e-08 2.166458402579977870409771e-19 -6.480960099352971832617487e-21 2.166458402579977870409771e-19 1.206246832769052560604811e-08 
1.206246832754287221234617e-08 9.071772495930309813082226e-20 -4.151557455857704423103985e-20 9.071772495930309813082226e-20 1.206246832769876763367159e-08 -1.400862420607288797217132e-19 -4.151557455857704423103985e-20 -1.400862420607288797217132e-19 1.206246832783158140718433e-08 
1.206246832768236464212466e-08 -1.813560405798011056048569e-19 -1.683167159859232320393665e-19 -1.813560405798011056048569e-19 1.206246832745240843183492e-08 9.117992505126417348521408e-20 -1.683167159859232320393665e-19 9.117992505126417348521408e-20 1.206246832793850442752416e-08 
  1.2062468327590134003825e-08 -4.548252598122822670280441e-20 -1.032066012452052790944902e-19 -4.548252598122822670280441e-20 1.206246832748899463032814e-08 -3.881607062951023841409701e-20 -1.032066012452052790944902e-19 -3.881607062951023841409701e-20 1.206246832799395530706726e-08 
1.206246832796692635337148e-08 1.467310873189439201624146e-19 1.639464607002770301192403e-19 1.467310873189439201624146e-19 1.206246832744081135964693e-08 4.125932951444460162663359e-20 1.639464607002770301192403e-19 4.125932951444460162663359e-20 1.206246832766560927163679e-08 
 1.20624683274664225257728e-08 -5.406617919769099488494501e-20 1.119497969223142124894216e-19 -5.406617919769099488494501e-20 1.206246832753729205193389e-08 4.993213729130410082285643e-20 1.119497969223142124894216e-19 4.993213729130410082285643e-20 1.206246832806961917205871e-08 
1.206246832751779209617356e-08 -7.20416410890808392875756e-20 -7.842227968976761423250009e-20 -7.20416410890808392875756e-20 1.206246832741129093794614e-08 6.464106294372203893741982e-20 -7.842227968976761423250009e-20 6.464106294372203893741982e-20  1.20624683281442904203151e-08 
1.206246832762205655802465e-08 -1.053604761627167940313959e-19 -6.254176579076768490073377e-20 -1.053604761627167940313959e-19 1.206246832757692558380375e-08 5.002788990955564934675151e-20 -6.254176579076768490073377e-20 5.002788990955564934675151e-20 1.206246832787426558115329e-08 
1.201671814753904965801822e-08 -5.806063437570956552689905e-20 1.081065090012397076550503e-19 -5.806063437570956552689905e-20 1.201671814733756335005133e-08 3.378495134880958583861038e-20 1.081065090012397076550503e-19 3.378495134880958583861038e-20  1.20167181475161235201607e-08 
1.201671814739777548120029e-08 6.520664768755517161011315e-20 5.763767043288220663756959e-20 6.520664768755517161011315e-20 1.201671814741878917748158e-08 6.831015179767170459988615e-20 5.763767043288220663756959e-20 6.831015179767170459988615e-20    1.201671814757614705413e-08 
1.201671814737799097530924e-08 -1.604151361924086569878123e-20 4.954377599371045432950431e-20 -1.604151361924086569878123e-20 1.201671814737735900932125e-08 -6.883073274630312411064351e-21 4.954377599371045432950431e-20 -6.883073274630312411064351e-21 1.201671814763751392941408e-08 
1.206246832742972217635504e-08 1.688503104889181567023135e-20 4.420784065728401105582757e-20 1.688503104889181567023135e-20 1.206246832793732817669311e-08 -1.033607153330815650631646e-19 4.420784065728401105582757e-20 -1.033607153330815650631646e-19 1.206246832770619240684987e-08 
1.206246832757324959316157e-08 -4.242526643723223641647968e-20 -1.539223499952355910876556e-20 -4.242526643723223641647968e-20 1.206246832749780741257428e-08 3.453737551350313363736529e-21 -1.539223499952355910876556e-20 3.453737551350313363736529e-21 1.206246832800249511971126e-08 
1.206246832748513500558997e-08 -4.166074475608010058797978e-20 3.382403563275271639624805e-20 -4.166074475608010058797978e-20 1.206246832786715182788534e-08 -1.573411262410084678910714e-20 3.382403563275271639624805e-20 -1.573411262410084678910714e-20 1.206246832772098570492476e-08 
1.206246832747909658711833e-08 -6.71521764882798927014107e-20 3.823568710753064923065793e-20 -6.71521764882798927014107e-20 1.206246832755020434129584e-08 -5.369848449071410294240725e-20 3.823568710753064923065793e-20 -5.369848449071410294240725e-20 1.206246832804405929113083e-08 
1.206246832787225222354234e-08 -1.158135575635494047587459e-19 1.702336925152306686421914e-19 -1.158135575635494047587459e-19 1.206246832746860959131239e-08 -3.369437507173502930821196e-20 1.702336925152306686421914e-19 -3.369437507173502930821196e-20 1.206246832773221385455956e-08 
1.206246832785757142203075e-08 -3.315199274408400906179878e-19 -2.50158442390124288517636e-19 -3.315199274408400906179878e-19 1.206246832742207902749505e-08 2.168228569090841349633995e-19 -2.50158442390124288517636e-19 2.168228569090841349633995e-19 1.206246832779366510226612e-08 
1.206246832742002265649225e-08 -1.088776481272922677049492e-19 4.882061334318596988474798e-20 -1.088776481272922677049492e-19  1.20624683275097816791216e-08 4.838324159429855650165972e-20 4.882061334318596988474798e-20 4.838324159429855650165972e-20 1.206246832814338217600252e-08 
1.201671814748885799280973e-08 4.951958096079327827001432e-20 4.907269663486150506866504e-20 4.951958096079327827001432e-20 1.201671814734956574073947e-08 -1.15362744129708004675941e-20 4.907269663486150506866504e-20 -1.15362744129708004675941e-20 1.201671814755420526120142e-08 
1.201671814745541508064421e-08 2.752443488270199588134612e-20 6.636325297905744255650209e-20 2.752443488270199588134612e-20 1.201671814738688316689419e-08 -4.670716687811298417545153e-20 6.636325297905744255650209e-20 -4.670716687811298417545153e-20 1.201671814755036548879794e-08 
1.201671814738605433192041e-08 -8.113152884042606040673751e-20 3.574909171331675005259254e-20 -8.113152884042606040673751e-20 1.201671814744801015980063e-08 -2.807187335184724650942196e-20 3.574909171331675005259254e-20 -2.807187335184724650942196e-20 1.201671814755874482840311e-08 
1.201671814738507660443637e-08 -2.868414210150134068151584e-20 4.715405120404475737680081e-20 -2.868414210150134068151584e-20 1.201671814738405751792171e-08 2.347124988119216027447622e-21 4.715405120404475737680081e-20 2.347124988119216027447622e-21 1.201671814762346013080681e-08 
1.206246832743596738997982e-08 -1.598485174728098330305254e-19 -7.823308797404025143398809e-20 -1.598485174728098330305254e-19 1.206246832750321055633548e-08 1.815931312228741171621669e-19 -7.823308797404025143398809e-20 1.815931312228741171621669e-19 1.206246832813409790080722e-08 
1.206246832765195748280721e-08 -2.043864031945025021286266e-19 1.475628432742601317716126e-19 -2.043864031945025021286266e-19 1.206246832762981385780917e-08 -1.318964043640237795591559e-19 1.475628432742601317716126e-19 -1.318964043640237795591559e-19 1.206246832779143502333468e-08 
1.201671814735876895223474e-08 1.000268155729748715838251e-21 -1.08185918340044798311838e-20 1.000268155729748715838251e-21 1.201671814737198895278456e-08 -4.311609149568472593557151e-20 -1.08185918340044798311838e-20 -4.311609149568472593557151e-20  1.20167181476619356098191e-08 
1.201671814738269432427222e-08 -9.643685171449473147488318e-21 4.331407200542046465312901e-20 -9.643685171449473147488318e-21 1.201671814739329877972515e-08 -1.462951631361284745777573e-20 4.331407200542046465312901e-20 -1.462951631361284745777573e-20 1.201671814761687908185333e-08 
!Field "H_trace" Scalar 1
3.605015444239257440083019e-08
3.618740498307340157857563e-08
3.618740498307315011566941e-08
 3.60501544423927266020629e-08
 3.60501544423927596892874e-08
3.605015444239266042761389e-08
3.618740498307329569945722e-08
 3.60501544423927530718425e-08
3.618740498307324937734292e-08
3.605015444239270013228329e-08
3.618740498307324937734292e-08
 3.60501544423928192462915e-08
3.618740498307333540412662e-08
3.618740498307315673311431e-08
3.618740498307340157857563e-08
3.605015444239261410549959e-08
3.605015444239262734038939e-08
3.605015444239302438708342e-08
3.618740498307313026333471e-08
  3.6050154442392719984618e-08
3.605015444239266042761389e-08
3.605015444239261410549959e-08
3.618740498307320967267352e-08
3.618740498307318982033881e-08
 3.60501544423928457160711e-08
3.605015444239267366250369e-08
3.618740498307340819602053e-08
3.605015444239268027994859e-08
 3.60501544423927464543976e-08
 3.60501544423927398369527e-08
3.618740498307329569945722e-08
 3.60501544423928324811813e-08
3.605015444239262734038939e-08
3.618740498307334202157152e-08
3.605015444239293174285481e-08
3.618740498307328908201232e-08
3.605015444239293174285481e-08
3.605015444239265381016899e-08
3.618740498307332216923682e-08
3.618740498307329569945722e-08
3.605015444239269351483839e-08
3.618740498307329569945722e-08
3.605015444239269351483839e-08
3.618740498307344128324503e-08
3.618740498307330231690212e-08
 3.60501544423927133671731e-08
3.618740498307325599478782e-08
 3.60501544423927927765119e-08
 3.60501544423928258637364e-08
3.605015444239303762197322e-08
3.618740498307326922967762e-08
3.618740498307324275989802e-08
3.618740498307333540412662e-08
 3.60501544423927266020629e-08
3.605015444239261410549959e-08
3.605015444239287880329561e-08
 3.60501544423928457160711e-08
3.605015444239266042761389e-08
3.605015444239286556840581e-08
3.618740498307321629011842e-08
3.605015444239269351483839e-08
3.618740498307329569945722e-08
 3.60501544423927596892874e-08
3.618740498307342143091033e-08
3.618740498307313688077961e-08
3.618740498307309717611021e-08
3.618740498307327584712252e-08
3.618740498307323614245312e-08
3.618740498307307070633061e-08
3.618740498307324937734292e-08
3.618740498307350084024913e-08
3.618740498307337510879603e-08
 3.60501544423927464543976e-08
3.618740498307332216923682e-08
3.618740498307322290756332e-08
3.618740498307321629011842e-08
3.618740498307327584712252e-08
3.618740498307308394122041e-08
3.618740498307334863901642e-08
3.618740498307333540412662e-08
3.618740498307337510879603e-08
3.618740498307324937734292e-08
 3.60501544423927398369527e-08
 3.60501544423927133671731e-08
3.605015444239286556840581e-08
3.618740498307324275989802e-08
3.618740498307355377980834e-08
3.618740498307327584712252e-08
3.618740498307336187390623e-08
3.618740498307307070633061e-08
3.618740498307331555179192e-08
3.618740498307318982033881e-08
3.605015444239262734038939e-08
3.605015444239266042761389e-08
 3.60501544423928126288466e-08
3.605015444239259425316489e-08
3.618740498307327584712252e-08
3.618740498307320967267352e-08
3.605015444239269351483839e-08
3.605015444239287218585071e-08
!Field "H_determinant" Scalar 1
1.735232306249560258231313e-24
1.755127043842946660539741e-24
1.755127043842909558999293e-24
1.735232306249582298750391e-24
1.735232306249586706854206e-24
1.735232306249573115200775e-24
1.755127043842930864834401e-24
1.735232306249585972170237e-24
1.755127043842923517994709e-24
1.735232306249578625330544e-24
1.755127043842923885336693e-24
1.735232306249595890403822e-24
 1.75512704384293710964814e-24
1.755127043842910661025247e-24
1.755127043842945925855771e-24
1.735232306249566135703067e-24
1.735232306249568339754975e-24
1.735232306249626012446562e-24
1.755127043842906620263416e-24
1.735232306249581931408406e-24
1.735232306249573115200775e-24
1.735232306249566870387036e-24
1.755127043842917640522955e-24
1.755127043842915069129062e-24
1.735232306249599931165653e-24
1.735232306249574584568713e-24
1.755127043842946660539741e-24
1.735232306249576421278637e-24
1.735232306249585604828252e-24
1.735232306249584502802299e-24
1.755127043842930130150432e-24
1.735232306249597359771761e-24
1.735232306249568339754975e-24
1.755127043842937476990125e-24
1.735232306249612420793131e-24
1.755127043842929395466463e-24
1.735232306249611686109161e-24
1.735232306249571278490852e-24
1.755127043842934170912263e-24
1.755127043842930497492417e-24
 1.73523230624957752330459e-24
1.755127043842930497492417e-24
1.735232306249577155962606e-24
 1.75512704384295217066951e-24
1.755127043842931232176386e-24
1.735232306249580462040468e-24
1.755127043842925354704632e-24
1.735232306249592216983976e-24
1.735232306249597359771761e-24
1.735232306249627849156485e-24
1.755127043842926456730586e-24
1.755127043842923150652724e-24
1.755127043842936742306156e-24
1.735232306249582298750391e-24
1.735232306249566503045052e-24
1.735232306249604339269469e-24
1.735232306249599563823668e-24
 1.73523230624957274785879e-24
1.735232306249602135217561e-24
1.755127043842919109890893e-24
1.735232306249577155962606e-24
1.755127043842930130150432e-24
1.735232306249587074196191e-24
1.755127043842948497249664e-24
  1.7551270438429069876054e-24
1.755127043842902579501585e-24
 1.75512704384292755875654e-24
 1.75512704384292204862677e-24
1.755127043842898171397769e-24
1.755127043842923517994709e-24
1.755127043842960619535157e-24
1.755127043842942252435925e-24
1.735232306249584870144283e-24
1.755127043842934538254248e-24
1.755127043842920211916847e-24
1.755127043842919844574863e-24
1.755127043842927926098524e-24
1.755127043842899640765708e-24
1.755127043842937844332109e-24
1.755127043842936007622186e-24
 1.75512704384294188509394e-24
1.755127043842923517994709e-24
1.735232306249583768118329e-24
1.735232306249580462040468e-24
1.735232306249602502559545e-24
 1.75512704384292278331074e-24
1.755127043842967599032865e-24
1.755127043842927191414555e-24
1.755127043842940048384017e-24
1.755127043842898538739754e-24
1.755127043842933436228294e-24
1.755127043842914701787078e-24
1.735232306249568339754975e-24
 1.73523230624957348254276e-24
1.735232306249594421035884e-24
1.735232306249563564309174e-24
 1.75512704384292755875654e-24
1.755127043842917640522955e-24
 1.73523230624957752330459e-24
1.735232306249603604585499e-24
!Field "H_eigen_min" Scalar 1
1.201671814746418981258217e-08
1.206246832769113441097895e-08
1.206246832769105003855647e-08
1.201671814746424109778015e-08
 1.20167181474642510239475e-08
1.201671800125984779898957e-08
  1.2062468327691098015032e-08
1.201671814746424936958627e-08
1.206246832769108147141975e-08
1.201671800125986268824059e-08
1.206246818093008164716468e-08
 1.20167181474642708762822e-08
1.206246832769111290428302e-08
1.206246832769105003855647e-08
1.206246812013973470641788e-08
1.201671800125983290973854e-08
1.201671814746420966491687e-08
1.201671814746434201381488e-08
1.206246832769104342111157e-08
1.201671814746424109778015e-08
1.201671814746422124544545e-08
 1.20167181474642047018332e-08
1.206246832769106823652995e-08
1.206246818093006179482998e-08
1.201671814746428245681078e-08
 1.20167181474642245541679e-08
1.206246832769113441097895e-08
1.201671814746422786289035e-08
1.201671814746424771522505e-08
1.201671789423084577035736e-08
1.206246832769109636067077e-08
1.201671800125990735599367e-08
1.201671814746420966491687e-08
1.206246832769111290428302e-08
1.201671800125994044321817e-08
1.206246832769109470630955e-08
1.201671814746430892659038e-08
1.201671814746421628236177e-08
1.206246832769110628683812e-08
  1.2062468327691098015032e-08
1.201671814746422951725157e-08
  1.2062468327691098015032e-08
1.201671814746422951725157e-08
1.206246832769114764586875e-08
  1.2062468327691098015032e-08
1.201671800125986599696304e-08
1.206246818093008330152591e-08
1.201671814746426260447608e-08
1.201671814746427583936588e-08
1.201671814746434532253733e-08
1.206246832769108808886465e-08
1.206246832769107981705852e-08
 1.20624683276911112499218e-08
1.201671814746424109778015e-08
1.201671814746420635619442e-08
1.201671814746429238297813e-08
1.201671814746428080244955e-08
1.201671814746421959108422e-08
1.201671814746428741989445e-08
1.206246832769107319961362e-08
1.201671814746422951725157e-08
1.206246832769109636067077e-08
1.201671814746425267830872e-08
1.206246832769113937406263e-08
1.206246832769104342111157e-08
1.206246832769103349494422e-08
 1.20624683276910913975871e-08
  1.2062468073493567435397e-08
1.206246832769102191441564e-08
1.206246832769108312578097e-08
1.206246832769116584384223e-08
1.206246832769112613917283e-08
1.201671814746424606086382e-08
1.206246832769110794119935e-08
1.206246832769107319961362e-08
1.206246818093007172099733e-08
 1.20624683276910913975871e-08
1.206246832769102687749932e-08
1.206246832769111621300547e-08
1.206246818093010977130551e-08
1.206246818093012300619531e-08
1.206246818093008164716468e-08
1.201671789423084577035736e-08
1.201671814746423613469647e-08
1.201671814746428741989445e-08
1.206246832769108147141975e-08
 1.20624683276911840418157e-08
 1.20624683276910913975871e-08
 1.20624683276911178673667e-08
1.206246818093002374452181e-08
 1.20624683276911046324769e-08
1.206246818093006179482998e-08
 1.20167181474642113192781e-08
1.201671814746421959108422e-08
1.201671814746426922192098e-08
1.201671800125982629229364e-08
 1.20624680734935806702868e-08
1.206246832769106989089117e-08
1.201671800125985937951814e-08
 1.20167181474642907286169e-08
!Field "H_eigen_max" Scalar 1
1.201671814746418981258217e-08
1.206246832769113441097895e-08
1.206246832769105003855647e-08
1.201671814746424109778015e-08
 1.20167181474642510239475e-08
1.201671843987296482963476e-08
  1.2062468327691098015032e-08
1.201671814746424936958627e-08
1.206246832769108147141975e-08
1.201671843987297806452456e-08
1.206246862121308773737477e-08
 1.20167181474642708762822e-08
1.206246832769111290428302e-08
1.206246832769105003855647e-08
1.206246874279393547446232e-08
1.201671843987294663166128e-08
1.201671814746420966491687e-08
1.201671814746434201381488e-08
1.206246832769104342111157e-08
1.201671814746424109778015e-08
1.201671814746422124544545e-08
 1.20167181474642047018332e-08
1.206246832769106823652995e-08
 1.20624686212130695394013e-08
1.201671814746428245681078e-08
 1.20167181474642245541679e-08
1.206246832769113441097895e-08
1.201671814746422786289035e-08
1.201671814746424771522505e-08
1.201671840069764635137029e-08
1.206246832769109636067077e-08
1.201671843987302273227763e-08
1.201671814746420966491687e-08
1.206246832769111290428302e-08
1.201671843987305416514091e-08
1.206246832769109470630955e-08
1.201671814746430892659038e-08
1.201671814746421628236177e-08
1.206246832769110628683812e-08
  1.2062468327691098015032e-08
1.201671814746422951725157e-08
  1.2062468327691098015032e-08
1.201671814746422951725157e-08
1.206246832769114764586875e-08
  1.2062468327691098015032e-08
1.201671843987298302760823e-08
1.206246862121309104609722e-08
1.201671814746426260447608e-08
1.201671814746427583936588e-08
1.201671814746434532253733e-08
1.206246832769108808886465e-08
1.206246832769107981705852e-08
 1.20624683276911112499218e-08
1.201671814746424109778015e-08
1.201671814746420635619442e-08
1.201671814746429238297813e-08
1.201671814746428080244955e-08
1.201671814746421959108422e-08
1.201671814746428741989445e-08
1.206246832769107319961362e-08
1.201671814746422951725157e-08
1.206246832769109636067077e-08
1.201671814746425267830872e-08
1.206246832769113937406263e-08
1.206246832769104342111157e-08
1.206246832769103349494422e-08
 1.20624683276910913975871e-08
1.206246858188859219872004e-08
1.206246832769102191441564e-08
1.206246832769108312578097e-08
1.206246832769116584384223e-08
1.206246832769112613917283e-08
1.201671814746424606086382e-08
1.206246832769110794119935e-08
1.206246832769107319961362e-08
1.206246862121307946556865e-08
 1.20624683276910913975871e-08
1.206246832769102687749932e-08
1.206246832769111621300547e-08
1.206246862121311751587683e-08
1.206246862121313075076663e-08
  1.2062468621213089391736e-08
1.201671840069764635137029e-08
1.201671814746423613469647e-08
1.201671814746428741989445e-08
1.206246832769108147141975e-08
 1.20624683276911840418157e-08
 1.20624683276910913975871e-08
 1.20624683276911178673667e-08
1.206246862121302983473189e-08
 1.20624683276911046324769e-08
1.206246862121306788504007e-08
 1.20167181474642113192781e-08
1.201671814746421959108422e-08
1.201671814746426922192098e-08
1.201671843987294001421638e-08
1.206246858188860543360984e-08
1.206246832769106989089117e-08
1.201671843987297475580211e-08
 1.20167181474642907286169e-08
!Field "work" Scalar 1
0.0001859999999999997777073296
0.0001529999999999997616247083
0.0001589999999999997719411088
0.0001539999999999997588265993
0.0001529999999999997616247083
0.0001499999999999997700190352
0.0001609999999999997663448909
0.0001519999999999997644228172
0.0001639999999999997850556183
0.0001489999999999997728171441
 0.000145999999999999781211471
0.0001519999999999997644228172
0.0001539999999999997588265993
0.0001479999999999997756152531
0.0001499999999999997700190352
0.0001479999999999997756152531
0.0001589999999999997719411088
0.0001669999999999997766612914
0.0001509999999999997672209262
0.0001539999999999997588265993
0.0001549999999999997560284903
0.0001539999999999997588265993
0.0001529999999999997887297626
0.0001479999999999997756152531
  0.00014499999999999978400958
0.0001469999999999997784133621
0.0001489999999999997728171441
0.0001519999999999997644228172
0.0001479999999999997756152531
0.0001519999999999997915278716
0.0001539999999999997588265993
0.0001569999999999997504322724
0.0001689999999999997710650734
0.0001509999999999997672209262
0.0001509999999999997943259805
0.0001509999999999997672209262
0.0001539999999999997588265993
0.0001599999999999997691429998
0.0001409999999999997952020159
0.0001479999999999997756152531
0.0001519999999999997644228172
0.0001509999999999997672209262
0.0001499999999999997700190352
0.0001469999999999997784133621
 0.000145999999999999781211471
0.0001679999999999997467581281
0.0001519999999999997644228172
0.0001499999999999997700190352
0.0001519999999999997644228172
0.0001559999999999997532303814
0.0001529999999999997616247083
0.0001509999999999997672209262
0.0001469999999999997784133621
 0.000145999999999999781211471
0.0001469999999999997784133621
0.0001519999999999997644228172
0.0001539999999999997588265993
0.0001659999999999997794594003
0.0001489999999999997728171441
0.0001489999999999997728171441
0.0001529999999999997616247083
0.0001679999999999997738631824
0.0001489999999999997728171441
0.0001499999999999997700190352
0.0001519999999999997644228172
0.0001499999999999997700190352
0.0001519999999999997644228172
0.0001469999999999997784133621
 0.000145999999999999781211471
0.0001469999999999997784133621
 0.000145999999999999781211471
0.0001499999999999997700190352
0.0001539999999999997588265993
0.0001569999999999997775373267
0.0001559999999999997532303814
0.0001529999999999997616247083
0.0001579999999999997476341634
0.0001529999999999997616247083
0.0001679999999999997738631824
0.0001529999999999997616247083
0.0001509999999999997672209262
0.0001669999999999997766612914
 0.000143999999999999786807689
0.0001499999999999997700190352
0.0001489999999999997728171441
0.0001559999999999997803354357
0.0001479999999999997756152531
0.0001499999999999997700190352
0.0001509999999999997672209262
0.0001519999999999997644228172
0.0001549999999999997560284903
0.0001529999999999997616247083
0.0001519999999999997644228172
0.0001649999999999997822575093
0.0001509999999999997672209262
0.0001539999999999997588265993
0.0001529999999999997616247083
0.0001519999999999997644228172
0.0001469999999999997784133621
0.0001469999999999997784133621
!Field "H_inverse" SymTensor 3 3
     83217396.6078859269618988 -0.0004981591417017882956336239 -0.0004361011974715937010438349 -0.0004981591417017882956336239     83217396.60799954831600189  2.73499473605050716991556e-05 -0.0004361011974715937010438349  2.73499473605050716991556e-05     83217396.60709628462791443 
    82901772.08086104691028595 0.0008668182392440044840842273 -0.0005335157096882746493790584 0.0008668182392440044840842273     82901772.07599884271621704  0.002255428719504753379970774 -0.0005335157096882746493790584  0.002255428719504753379970774      82901772.0770544707775116 
    82901772.07833786308765411 -0.001358258084335799403125078 -0.0006979889213637978373494519 -0.001358258084335799403125078      82901772.0770760178565979 -0.0001005983397386354732602753 -0.0006979889213637978373494519 -0.0001005983397386354732602753     82901772.07850223779678345 
    83217396.60865224897861481 0.0002174820612455083824587215 7.677833949687404302159727e-05 0.0002174820612455083824587215     83217396.60843861103057861 0.0004460176657098001602730353 7.677833949687404302159727e-05 0.0004460176657098001602730353     83217396.60588982701301575 
    83217396.60812371969223022 6.277112224307004938270854e-05 -0.0004469678536936523278837174 6.277112224307004938270854e-05     83217396.60817337036132812 0.0001012268839135395804944284 -0.0004469678536936523278837174 0.0001012268839135395804944284     83217396.60668341815471649 
    83217396.60816812515258789 -0.0003472002637621400414694173 -3.610642725785319140157856e-05 -0.0003472002637621400414694173     83217396.60806766152381897 0.0001390152942674304469006241 -3.610642725785319140157856e-05 0.0001390152942674304469006241     83217396.60674537718296051 
    82901772.07883095741271973 0.0005958357430457618180916213 0.0003356362086390876652876314 0.0005958357430457618180916213     82901772.07872167229652405 -0.0006986064509266897044892364 0.0003356362086390876652876314 -0.0006986064509266897044892364     82901772.07636247575283051 
    83217396.60810528695583344 5.651577770107883897689194e-05 -0.0004683288242030791644933407 5.651577770107883897689194e-05     83217396.60817252099514008 0.0001123377105224229532227584 -0.0004683288242030791644933407 0.0001123377105224229532227584     83217396.60670273005962372 
    82901772.07866045832633972 0.0004799363136712915035332616 0.0003928873829633342971631715 0.0004799363136712915035332616      82901772.0791100412607193 -0.0004145094456620629971149716 0.0003928873829633342971631715 -0.0004145094456620629971149716     82901772.07614494860172272 
    83217396.60842834413051605 0.0004040597417158412136065082 4.127714689788128281172034e-06 0.0004040597417158412136065082     83217396.60832720994949341 2.147441844330911435261011e-05 4.127714689788128281172034e-06 2.147441844330911435261011e-05     83217396.60622534155845642 
    82901772.07847622036933899 0.0009276104376183306153558217 7.327567604069695306016896e-05 0.0009276104376183306153558217     82901772.07810743153095245 -0.0002096750976812638623310997 7.327567604069695306016896e-05 -0.0002096750976812638623310997      82901772.0773317813873291 
    83217396.60829968750476837 0.0002053150724089704975972026 -0.0001607841403065430468943831 0.0002053150724089704975972026     83217396.60823886096477509 0.0002188425413928601925318829 -0.0001607841403065430468943831 0.0002188425413928601925318829     83217396.60644151270389557 
    82901772.07749137282371521  0.001563650269753058411406621 -0.001304666963023168270094376  0.001563650269753058411406621     82901772.07937522232532501 0.0009762581244523382221350838 -0.001304666963023168270094376 0.0009762581244523382221350838     82901772.07704819738864899 
    82901772.07958625257015228  0.000184383388570374972571797 0.0001052815092583400847928501  0.000184383388570374972571797     82901772.08006297051906586 0.0001295980688239708837877079 0.0001052815092583400847928501 0.0001295980688239708837877079     82901772.07426685094833374 
    82901772.07860876619815826  0.001712761278392490628397216 -2.952629918856345195288249e-05  0.001712761278392490628397216     82901772.07759580016136169 -0.0005733886494498314579174036 -2.952629918856345195288249e-05 -0.0005733886494498314579174036     82901772.07770980894565582 
    83217396.60732182860374451 -0.0003848268485808281689879162 -0.0004514409692321202363304855 -0.0003848268485808281689879162     83217396.60848855972290039 0.0001434518916587454071768365 -0.0004514409692321202363304855 0.0001434518916587454071768365     83217396.60717108845710754 
     83217396.6076444685459137                              0                              0                              0     83217396.60846564173698425                              0                              0                              0     83217396.60687126219272614 
    83217396.60836827754974365 -0.0002703202462745221516804417 -0.0001658654441805448419983149 -0.0002703202462745221516804417     83217396.60776445269584656 0.0002715439623664004493118485 -0.0001658654441805448419983149 0.0002715439623664004493118485     83217396.60684587061405182 
    82901772.07933114469051361 -0.0003584101878543610058582003 -0.0001292519964415549322319515 -0.0003584101878543610058582003     82901772.07680514454841614 0.0002164794706332128198644077 -0.0001292519964415549322319515 0.0002164794706332128198644077     82901772.07777997851371765 
    83217396.60848341882228851 0.0003355831953287259335552695 -0.0002071130543335367819521298 0.0003355831953287259335552695      83217396.6083768755197525 0.0003789005254161107328486624 -0.0002071130543335367819521298 0.0003789005254161107328486624     83217396.60612042248249054 
    83217396.60830837488174438 0.0006366474289250997073766336 0.0001031143711151298131495704 0.0006366474289250997073766336     83217396.60811397433280945 -0.000330684750721817915294215 0.0001031143711151298131495704 -0.000330684750721817915294215     83217396.60655881464481354 
    83217396.60826894640922546 0.0002085974097928802750180621 -0.0003307413180557554626022576 0.0002085974097928802750180621     83217396.60825009644031525 -7.096121277309768457606381e-05 -0.0003307413180557554626022576 -7.096121277309768457606381e-05     83217396.60646238923072815 
    82901772.07692234218120575 0.0003158653134455427133851779 -0.0005719491091186899769244212 0.0003158653134455427133851779     82901772.07927447557449341 -8.444734751103412232538931e-05 -0.0005719491091186899769244212 -8.444734751103412232538931e-05     82901772.07771891355514526 
    82901772.07978911697864532 -0.0004985844278086728684207252 -0.0004473017585952511693606071 -0.0004985844278086728684207252      82901772.0758003443479538 -0.0006128366378825313674771902 -0.0004473017585952511693606071 -0.0006128366378825313674771902     82901772.07832640409469604 
    83217396.60857079923152924 0.0003817707805298085638884276 -0.0005391138905952244392977279 0.0003817707805298085638884276     83217396.60825362801551819 0.0004049726954898316580271078 -0.0005391138905952244392977279 0.0004049726954898316580271078     83217396.60615544021129608 
    83217396.60813350975513458 3.049766880985738291766525e-05 -0.0004365193661066805747711372 3.049766880985738291766525e-05     83217396.60831433534622192 0.0001250474593339683871458939 -0.0004365193661066805747711372 0.0001250474593339683871458939      83217396.6065332442522049 
    82901772.07876439392566681 0.0002889612054639645408876669 -0.000234619468620248465941594 0.0002889612054639645408876669     82901772.07905110716819763 0.0001353887410363041631823633 -0.000234619468620248465941594 0.0001353887410363041631823633     82901772.07609887421131134 
    83217396.60851305723190308 -2.962177020547271310223734e-05 -0.0002427354370768860223651908 -2.962177020547271310223734e-05     83217396.60741351544857025 -4.44833152922372994614135e-05 -0.0002427354370768860223651908 -4.44833152922372994614135e-05     83217396.60705441236495972 
    83217396.60723978281021118 0.0004109308825330586201728111 -8.006998542636700689958257e-05 0.0004109308825330586201728111     83217396.60850532352924347 0.0001776686835836845243172255 -8.006998542636700689958257e-05 0.0001776686835836845243172255     83217396.60723543167114258 
    83217396.60818788409233093 9.579498788821090300271005e-05 -0.0002893956101195602507655802 9.579498788821090300271005e-05     83217396.60817034542560577 4.484643818602274876984268e-05 -0.0002893956101195602507655802 4.484643818602274876984268e-05      83217396.6066223531961441 
    82901772.07864393293857574 0.0004212219708763886133993937 -0.0003890531389680245235619671 0.0004212219708763886133993937     82901772.07940959930419922 0.0002552813270067438378499447 -0.0003890531389680245235619671 0.0002552813270067438378499447     82901772.07586164772510529 
    83217396.60849873721599579 0.0001691749911690613940480621 -0.0004583099619272111222012533 0.0001691749911690613940480621     83217396.60843849182128906 7.175315542947064730017193e-05 -0.0004583099619272111222012533 7.175315542947064730017193e-05      83217396.6060427725315094 
    83217396.60850369930267334 0.0002380639778557750861794073 -0.000116243720650484401077894 0.0002380639778557750861794073      83217396.6083921492099762 -0.0001613314650532550378198016 -0.000116243720650484401077894 -0.0001613314650532550378198016     83217396.60608549416065216 
    82901772.07776761054992676 -0.001214286286194752977063427 -0.0005186495200745468376127278 -0.001214286286194752977063427     82901772.07824802398681641 -9.345375702542475641367015e-05 -0.0005186495200745468376127278 -9.345375702542475641367015e-05     82901772.07789914309978485 
    83217396.60822699964046478 7.646184885020277321142357e-05 -0.0002413592039918836243059252 7.646184885020277321142357e-05     83217396.60817071795463562 0.0002595076512311508950756056 -0.0002413592039918836243059252 0.0002595076512311508950756056     83217396.60658150911331177 
    82901772.07699751853942871 -3.148441511787244831768739e-05 -0.0007079035044060377323410505 -3.148441511787244831768739e-05     82901772.07926908135414124 -7.221542963287704388394145e-05 -0.0007079035044060377323410505 -7.221542963287704388394145e-05      82901772.0776485800743103 
     83217396.6081443727016449 0.0001497101003680112397877661 -0.0002346288661525245311436499 0.0001497101003680112397877661      83217396.6082228422164917 0.0001799693215330584630633204 -0.0002346288661525245311436499 0.0001799693215330584630633204     83217396.60661210119724274 
    83217396.60851027071475983                             -0                             -0                             -0     83217396.60787773132324219 0.0004712560046598992320905641                             -0 0.0004712560046598992320905641     83217396.60659325122833252 
    82901772.07773977518081665  0.002251110631577695267435679 0.0009248034849601117568865249  0.002251110631577695267435679     82901772.07851362228393555 -0.0005852254620747861842827708 0.0009248034849601117568865249 -0.0005852254620747861842827708     82901772.07766157388687134 
    82901772.07856474816799164 -0.0006671650283865007777933664 -0.0009647695160575109384407111 -0.0006671650283865007777933664     82901772.07902386784553528 -0.0008854237161311397227500541 -0.0009647695160575109384407111 -0.0008854237161311397227500541     82901772.07632648944854736 
    83217396.60819973051548004 0.0005316240893324893947158305 -0.0003603131443164443920880446 0.0005316240893324893947158305     83217396.60792946815490723 0.0004983781610965463178958279 -0.0003603131443164443920880446 0.0004983781610965463178958279       83217396.606851726770401 
    82901772.08041539788246155 0.0005564275493982103739862288 -0.0004193629865531301511433204 0.0005564275493982103739862288     82901772.07900811731815338 -0.002252169456681263164099516 -0.0004193629865531301511433204 -0.002252169456681263164099516     82901772.07449162006378174 
    83217396.60798667371273041 -0.0001652682649980363087729995 -0.0003584349656635419452584135 -0.0001652682649980363087729995      83217396.6081211268901825 4.450918231730640397007456e-05 -0.0003584349656635419452584135 4.450918231730640397007456e-05     83217396.60687315464019775 
    82901772.07880426943302155 0.0002969684819799445012721006 -0.0002091234337769820768315743 0.0002969684819799445012721006     82901772.07965824007987976 2.394259530603881085835706e-05 -0.0002091234337769820768315743 2.394259530603881085835706e-05     82901772.07545159757137299 
    82901772.07725836336612701  0.001942303205096968963735971 -0.001028234359703555185136525  0.001942303205096968963735971     82901772.07871416211128235 9.302312073270250190881736e-05 -0.001028234359703555185136525 9.302312073270250190881736e-05     82901772.07794253528118134 
    83217396.60849820077419281 0.0005528303947317710640221855 -0.0004158386356729431828152532 0.0005528303947317710640221855      83217396.6079629510641098 0.0005090118350910205003226339 -0.0004158386356729431828152532 0.0005090118350910205003226339     83217396.60651962459087372 
    82901772.07827125489711761  0.001097090684274242737908378 -0.0005578587398913073449463473  0.001097090684274242737908378     82901772.07842786610126495 -3.256633547452053134129563e-05 -0.0005578587398913073449463473 -3.256633547452053134129563e-05      82901772.0772162526845932 
    83217396.60823579132556915 7.743566622459584268631932e-05 -0.0002896920515847880672581638 7.743566622459584268631932e-05      83217396.6081782728433609 3.256559864439972852741267e-05 -0.0002896920515847880672581638 3.256559864439972852741267e-05      83217396.6065661609172821 
    83217396.60860691964626312  0.000111112562345940188717093 0.0003718736454188664047361412  0.000111112562345940188717093      83217396.6086353212594986 0.0002778959726025138346136578 0.0003718736454188664047361412 0.0002778959726025138346136578     83217396.60573774576187134 
    83217396.60840624570846558                             -0                             -0                             -0     83217396.60835924744606018 0.0001974715462929992613235614                             -0 0.0001974715462929992613235614      83217396.6062130331993103 
    82901772.07585564255714417 -0.0007559869582660187770084548 0.0001030488715724808877847313 -0.0007559869582660187770084548     82901772.07992476224899292 3.479102308115569953299653e-05 0.0001030488715724808877847313 3.479102308115569953299653e-05      82901772.0781349241733551 
    82901772.07920356094837189  0.000303668215998518381277399 -0.0001464760262713385777482572  0.000303668215998518381277399     82901772.07782050967216492 -0.0005840078131457412729740653 -0.0001464760262713385777482572 -0.0005840078131457412729740653     82901772.07689142227172852 
    82901772.07992440462112427 0.0005055641464940433633598604 -0.0002828178876084393167378295 0.0005055641464940433633598604     82901772.07884253561496735 0.0005399847583914982275185568 -0.0002828178876084393167378295 0.0005399847583914982275185568     82901772.07514789700508118 
    83217396.60838395357131958 0.0007752617395641003524356383 -0.0003638917441540135593383565 0.0007752617395641003524356383      83217396.6075565367937088 0.0005505605409871532551421835 -0.0003638917441540135593383565 0.0005505605409871532551421835     83217396.60704021155834198 
    83217396.60831281542778015 -0.0004270819300904859648800038  0.000740427808764807719558998 -0.0004270819300904859648800038     83217396.60824243724346161 0.0007983651092159604846162924  0.000740427808764807719558998 0.0007983651092159604846162924     83217396.60642623901367188 
     83217396.6085212230682373 -5.820814340837771825578825e-05 -0.0002591442598206798882641555 -5.820814340837771825578825e-05     83217396.60842595994472504 -0.0005661946060907059510153294 -0.0002591442598206798882641555 -0.0005661946060907059510153294     83217396.60603244602680206 
    83217396.60810001194477081  3.32673199880515030302762e-05 -0.0003662330230954933879203295  3.32673199880515030302762e-05     83217396.60827341675758362 2.183069418367710354494764e-05 -0.0003662330230954933879203295 2.183069418367710354494764e-05     83217396.60660648345947266 
    83217396.60835522413253784 0.0002225630965990350624162525 -0.0003545941153732466146961122 0.0002225630965990350624162525     83217396.60833431780338287 0.0002227317245284510347381329 -0.0003545941153732466146961122 0.0002227317245284510347381329     83217396.60629165172576904 
    83217396.60808348655700684  4.24183391322014262934427e-05 -0.0003670950036302397800902497  4.24183391322014262934427e-05     83217396.60825757682323456  7.32777882563050196942922e-05 -0.0003670950036302397800902497  7.32777882563050196942922e-05     83217396.60663869976997375 
    82901772.07795199751853943 0.0009840678484016429205388787  0.001981256601316029770931681 0.0009840678484016429205388787     82901772.08076639473438263 -1.33838343613654363784167e-05  0.001981256601316029770931681 -1.33838343613654363784167e-05     82901772.07519726455211639 
    83217396.60809117555618286 0.0001423090883280696532925402 -0.0004608461833534793707263522 0.0001423090883280696532925402     83217396.60820247232913971 -1.573860726136594909130816e-05 -0.0004608461833534793707263522 -1.573860726136594909130816e-05     83217396.60668729245662689 
    82901772.07919564843177795 0.0008860789086338038272883111 -0.0005092480053183977544567496 0.0008860789086338038272883111     82901772.07728847861289978 0.0007092252593102173555128509 -0.0005092480053183977544567496 0.0007092252593102173555128509     82901772.07743103802204132 
    83217396.60811826586723328 0.0005242689039958247461045704 9.540868312579280910087909e-05 0.0005242689039958247461045704     83217396.60829786956310272 -0.0001582968782664287573334894 9.540868312579280910087909e-05 -0.0001582968782664287573334894     83217396.60656434297561646 
    82901772.07684582471847534 -0.0008345702619514740487269289 -0.0009371085967955963130782138 -0.0008345702619514740487269289     82901772.07920660078525543 -0.0002593467892813920683790785 -0.0009371085967955963130782138 -0.0002593467892813920683790785     82901772.07786186039447784 
    82901772.07729226350784302  0.001043799800323620078496001 -0.001283489082824859671763673  0.001043799800323620078496001     82901772.07951436936855316 0.0005051794340667325588362102 -0.001283489082824859671763673 0.0005051794340667325588362102     82901772.07710961997509003 
    82901772.07585608959197998 -0.0006046474424288844759164951  -0.00076456841646732522782548 -0.0006046474424288844759164951     82901772.07976582646369934 0.0001032887505573455542854169  -0.00076456841646732522782548 0.0001032887505573455542854169     82901772.07829450070858002 
    82901772.07952871918678284  0.001159920943420000372450773 -0.0007779039286387140310352617  0.001159920943420000372450773     82901772.07704414427280426  0.001107707360759368217864584 -0.0007779039286387140310352617  0.001107707360759368217864584     82901772.07734240591526031 
    82901772.07971121370792389   0.00018631911997152425432972  0.001137940017132848787365096   0.00018631911997152425432972     82901772.08022983372211456  0.001291761021222153802898158  0.001137940017132848787365096  0.001291761021222153802898158     82901772.07397447526454926 
     82901772.0786176323890686 0.0006586603172348785969689167 -0.0005876088846530464447626141 0.0006586603172348785969689167     82901772.07857999205589294 0.0003279956125208746036195362 -0.0005876088846530464447626141 0.0003279956125208746036195362      82901772.0767190009355545 
    82901772.07917216420173645 -0.0004897855195948596111407691 -0.000647432506706678871297167 -0.0004897855195948596111407691     82901772.07765170931816101 -0.000990640381228936970497978 -0.000647432506706678871297167 -0.000990640381228936970497978     82901772.07709160447120667 
    82901772.07972529530525208 0.0004344849997176091611038318 0.0002935276554813085782280613 0.0004344849997176091611038318     82901772.07972754538059235  0.001036184786534200506780135 0.0002935276554813085782280613  0.001036184786534200506780135     82901772.07446087896823883 
    82901772.07952864468097687 0.0004793962417814484752373594 -0.0009116598404555446713906641 0.0004793962417814484752373594     82901772.07914118468761444 -0.0001182146323308819814727408 -0.0009116598404555446713906641 -0.0001182146323308819814727408      82901772.0752447247505188 
    83217396.60836711525917053 0.0003403606287987803518876873 0.0002252110206001122015128518 0.0003403606287987803518876873     83217396.60852465033531189  5.34303519196272167228641e-05 0.0002252110206001122015128518  5.34303519196272167228641e-05     83217396.60608881711959839 
    82901772.07957898080348969  0.001353434389544084419723657 -5.195704848287799478522009e-05  0.001353434389544084419723657     82901772.07609118521213531 -0.0001750008829131361549804463 -5.195704848287799478522009e-05 -0.0001750008829131361549804463     82901772.07824476063251495 
    82901772.08000998198986053  0.001276167155803460120586101  4.45417191692299791134016e-05  0.001276167155803460120586101     82901772.07592998445034027 -0.001488942692519158164307647  4.45417191692299791134016e-05 -0.001488942692519158164307647     82901772.07797564566135406 
    82901772.07899041473865509 -0.0006234760542990357319592665 0.0002853242475882919308195762 -0.0006234760542990357319592665     82901772.07791900634765625 0.0009627712500392148799177594 0.0002853242475882919308195762 0.0009627712500392148799177594     82901772.07700622081756592 
    82901772.07803173363208771  0.001246406351741344200462214  0.001156790935828212870881138  0.001246406351741344200462214     82901772.07961215078830719 -0.0006266526186119381535907791  0.001156790935828212870881138 -0.0006266526186119381535907791     82901772.07627135515213013 
     82901772.0786655992269516  0.000312587929776576010140049 0.0007093084019627657723153225  0.000312587929776576010140049      82901772.0793607085943222 0.0002667713566474865655164805 0.0007093084019627657723153225 0.0002667713566474865655164805     82901772.07589027285575867 
    82901772.07607603073120117 -0.001008439303394564542926126 -0.001126755465665326512089695 -0.001008439303394564542926126     82901772.07969187200069427 -0.0002835631512960835941099258 -0.001126755465665326512089695 -0.0002835631512960835941099258     82901772.07814688980579376 
    82901772.07951584458351135 0.0003715808359772706875000237 -0.0007693977962390688256355542 0.0003715808359772706875000237     82901772.07902878522872925 -0.0003431687903835940007743477 -0.0007693977962390688256355542 -0.0003431687903835940007743477     82901772.07537025213241577 
    82901772.07916279137134552 0.0004951208614715354268051573  0.000538973100685242903322425 0.0004951208614715354268051573     82901772.07989473640918732 -0.0004442588798032650731356652  0.000538973100685242903322425 -0.0004442588798032650731356652     82901772.07485705614089966 
    82901772.07844622433185577 0.0007241113463425926733210702 0.0004298310322566681871726824 0.0007241113463425926733210702     82901772.07875639200210571 -0.0003438268697654434623289799 0.0004298310322566681871726824 -0.0003438268697654434623289799     82901772.07671286165714264 
    83217396.60714218020439148 0.0004020777369403056330891821 -0.000748652179816907390776104 0.0004020777369403056330891821     83217396.60853751003742218 -0.0002339653523802286887254415 -0.000748652179816907390776104 -0.0002339653523802286887254415     83217396.60730095207691193 
    83217396.60812051594257355 -0.0004515648445361582392909572 -0.0003991486544866603911052572 -0.0004515648445361582392909572     83217396.60797499120235443 -0.0004730570297696808958198833 -0.0003991486544866603911052572 -0.0004730570297696808958198833     83217396.60688526928424835 
    83217396.60825753211975098 0.0001110896489935663867566762 -0.0003430973420267054586202393 0.0001110896489935663867566762     83217396.60826189815998077 4.766621231652550650216907e-05 -0.0003430973420267054586202393 4.766621231652550650216907e-05     83217396.60646030306816101 
    82901772.07976807653903961 -0.0001160458172863700141829585 -0.0003038273950865394423814791 -0.0001160458172863700141829585     82901772.07627944648265839 0.0007103675824381549402941616 -0.0003038273950865394423814791 0.0007103675824381549402941616     82901772.07786796987056732 
    82901772.07878166437149048  0.000291576290446536384379228  0.000105786272180318315820971  0.000291576290446536384379228      82901772.0793001651763916 -2.373651523996910605121026e-05  0.000105786272180318315820971 -2.373651523996910605121026e-05     82901772.07583159208297729 
    82901772.07938723266124725 0.0002863219593657663247961154 -0.0002324625786898806942444573 0.0002863219593657663247961154     82901772.07676175236701965 0.0001081358958336901815574724 -0.0002324625786898806942444573 0.0001081358958336901815574724      82901772.0777662992477417 
    82901772.07942873239517212 0.0004615170194594379600265543 -0.0002627825525970157592887955 0.0004615170194594379600265543     82901772.07894003391265869 0.0003690537791395699651619822 -0.0002627825525970157592887955 0.0003690537791395699651619822     82901772.07554592192173004 
    82901772.07672670483589172 0.0007959522787409204803987794 -0.001169965747740424723624675 0.0007959522787409204803987794     82901772.07950082421302795 0.0002315714600469212351447484 -0.001169965747740424723624675 0.0002315714600469212351447484     82901772.07768914103507996 
    82901772.07682758569717407  0.002278438269618055997400852  0.001719264880956545204701569  0.002278438269618055997400852     82901772.07982060313224792  -0.00149015927554275854662047  0.001719264880956545204701569  -0.00149015927554275854662047     82901772.07726681232452393 
    82901772.07983472943305969 0.0007482838275370503645922415 -0.0003355296155072845639896761 0.0007482838275370503645922415     82901772.07921783626079559 -0.0003325236890183133121358383 -0.0003355296155072845639896761 -0.0003325236890183133121358383     82901772.07486329972743988 
    83217396.60748976469039917 -0.0003429297881604942356721655 -0.0003398350538243606329229241 -0.0003429297881604942356721655      83217396.6084543764591217 7.989025884079498486881055e-05 -0.0003398350538243606329229241 7.989025884079498486881055e-05     83217396.60703721642494202 
    83217396.60772135853767395 -0.0001906104300662794022881014 -0.0004595744924309023439999711 -0.0001906104300662794022881014      83217396.6081959456205368 0.0003234534406838953215015953 -0.0004595744924309023439999711 0.0003234534406838953215015953     83217396.60706381499767303 
    83217396.60820168256759644 0.0005618467979437768771919237 -0.0002475672897494612099446309 0.0005618467979437768771919237     83217396.60777264833450317 0.0001944015154169472111254924 -0.0002475672897494612099446309 0.0001944015154169472111254924       83217396.607005774974823 
    83217396.60820844769477844 0.0001986415592303168373145006 -0.0003265481750112681912263934 0.0001986415592303168373145006     83217396.60821551084518433 -1.62541576356573965725285e-05 -0.0003265481750112681912263934 -1.62541576356573965725285e-05     83217396.60655762255191803 
    82901772.07972516119480133   0.00109859151567680518417347 0.0005376728420492955231799193   0.00109859151567680518417347     82901772.07926301658153534 -0.001248035805457834964207753 0.0005376728420492955231799193 -0.001248035805457834964207753     82901772.07492710649967194 
    82901772.07824070751667023  0.001404687212697342110420684 -0.001014155715706191885489007  0.001404687212697342110420684     82901772.07839290797710419 0.0009064849212616001451064962 -0.001014155715706191885489007 0.0009064849212616001451064962     82901772.07728211581707001 
    83217396.60839065909385681 -6.926992112657640717160532e-06 7.492021002169521961839421e-05 -6.926992112657640717160532e-06     83217396.60829910635948181 0.0002985847585094723670960659 7.492021002169521961839421e-05 0.0002985847585094723670960659     83217396.60629118978977203 
    83217396.60822495818138123 6.678382265685959954561179e-05 -0.0002999558002869645969082346 6.678382265685959954561179e-05     83217396.60815152525901794 0.0001013113768915257259344009 -0.0002999558002869645969082346 0.0001013113768915257259344009     83217396.60660319030284882 
!Field "H_inverse_trace" Scalar 1
    249652189.8229817450046539
    248705316.2339143455028534
    248705316.2339161038398743
     249652189.822980672121048
     249652189.822980523109436
    249652189.8229811787605286
    248705316.2339150905609131
     249652189.822980523109436
    248705316.2339154481887817
    249652189.8229809105396271
    248705316.2339154481887817
    249652189.8229800462722778
    248705316.2339147925376892
    248705316.2339160740375519
    248705316.2339143753051758
    249652189.8229814767837524
    249652189.8229813575744629
    249652189.8229786157608032
    248705316.2339162528514862
    249652189.8229807019233704
    249652189.8229811787605286
    249652189.8229814469814301
    248705316.2339157462120056
    248705316.2339158654212952
    249652189.8229798674583435
     249652189.822981059551239
    248705316.2339143753051758
    249652189.8229809999465942
     249652189.822980523109436
    249652189.8229805827140808
    248705316.2339151501655579
    249652189.8229800164699554
    249652189.8229813575744629
    248705316.2339147925376892
     249652189.822979211807251
    248705316.2339151799678802
    249652189.8229793310165405
    249652189.8229812383651733
    248705316.2339149713516235
    248705316.2339150905609131
    249652189.8229809105396271
    248705316.2339151501655579
    249652189.8229809403419495
    248705316.2339141368865967
    248705316.2339150905609131
    249652189.8229807615280151
     248705316.233915388584137
    249652189.8229802250862122
    249652189.8229799866676331
    249652189.8229785263538361
    248705316.2339153289794922
    248705316.2339155077934265
    248705316.2339148223400116
    249652189.8229807019233704
    249652189.8229814767837524
    249652189.8229796290397644
    249652189.8229799270629883
    249652189.8229811787605286
    249652189.8229797780513763
    248705316.2339156866073608
    249652189.8229809403419495
    248705316.2339151501655579
    249652189.8229804635047913
    248705316.2339142560958862
    248705316.2339162826538086
    248705316.2339164018630981
    248705316.2339152693748474
    248705316.2339155077934265
    248705316.2339166402816772
    248705316.2339154779911041
    248705316.2339137196540833
    248705316.2339145541191101
    249652189.8229805827140808
    248705316.2339149117469788
    248705316.2339156270027161
    248705316.2339156270027161
     248705316.233915239572525
    248705316.2339165806770325
    248705316.2339147925376892
    248705316.2339148819446564
    248705316.2339145839214325
    248705316.2339154481887817
    249652189.8229806423187256
    249652189.8229807615280151
    249652189.8229797184467316
    248705316.2339155077934265
    248705316.2339134216308594
    248705316.2339152693748474
    248705316.2339146733283997
    248705316.2339166700839996
    248705316.2339150011539459
    248705316.2339158654212952
    249652189.8229813575744629
    249652189.8229811191558838
    249652189.8229801058769226
     249652189.822981595993042
    248705316.2339152693748474
    248705316.2339157462120056
    249652189.8229809403419495
    249652189.8229796886444092
!Field "H_inverse_determinant" Scalar 1
      576291714024934897352704
      569759325120103742177280
      569759325120115754663936
      576291714024927448268800
      576291714024926307418112
      576291714024930803712000
      569759325120108775342080
      576291714024926441635840
      569759325120111191261184
      576291714024928924663808
      569759325120111057043456
      576291714024923220410368
      569759325120106694967296
      569759325120115419119616
      569759325120103742177280
      576291714024933018304512
      576291714024932280107008
      576291714024913019863040
      569759325120116828405760
      576291714024927716704256
      576291714024930870820864
      576291714024932615651328
      569759325120113137418240
      569759325120114009833472
      576291714024921878233088
      576291714024930266841088
      569759325120103809286144
      576291714024929528643584
      576291714024926441635840
      576291714024926777180160
      569759325120109312212992
      576291714024922817757184
      576291714024932078780416
      569759325120106627858432
      576291714024917381939200
      569759325120109312212992
      576291714024918053027840
      576291714024931407691776
      569759325120107970035712
      569759325120108842450944
      576291714024929125990400
      569759325120109043777536
      576291714024929394425856
      569759325120101997346816
      569759325120108506906624
      576291714024928119357440
      569759325120110654390272
      576291714024924294152192
      576291714024922683539456
      576291714024912550100992
      569759325120110385954816
      569759325120111526805504
      569759325120107030511616
      576291714024927649595392
      576291714024933085413376
      576291714024920200511488
      576291714024922146668544
      576291714024931005038592
      576291714024921072926720
      569759325120112600547328
      576291714024929327316992
      569759325120109177995264
      576291714024926106091520
      569759325120103205306368
      569759325120116761296896
      569759325120117835038720
      569759325120109983301632
      569759325120111661023232
      569759325120119311433728
      569759325120111392587776
      569759325120099312992256
      569759325120105017245696
      576291714024926777180160
      569759325120107634491392
      569759325120112332111872
      569759325120112533438464
      569759325120109714866176
      569759325120118975889408
      569759325120106627858432
      569759325120107298947072
      569759325120105218572288
      569759325120111325478912
      576291714024927246942208
      576291714024928119357440
      576291714024920938708992
      569759325120111459696640
      569759325120097232617472
      569759325120110117519360
      569759325120105889660928
      569759325120119579869184
      569759325120108037144576
      569759325120114076942336
      576291714024932145889280
      576291714024930468167680
      576291714024923488845824
      576291714024933756502016
      569759325120110050410496
      569759325120113070309376
      576291714024929327316992
      576291714024920536055808
!Field "H_inverse_eigen_min" Scalar 1
    83217396.60766057670116425
     82901772.0779714435338974
    82901772.07797203958034515
    83217396.60766021907329559
    83217395.59517514705657959
    83217396.60766038298606873
     82901772.0779716968536377
    83217394.85398468375205994
    82901772.07797181606292725
    83217396.60766029357910156
    82901771.06932692229747772
    83217396.60766001045703888
     82901770.3309473842382431
    82901772.07797202467918396
    82901772.07797145843505859
    83217396.60766048729419708
    83217395.59517543017864227
    83217396.60765953361988068
    82901772.07797208428382874
    83217396.60766023397445679
    83217396.60766036808490753
    83217396.60766047239303589
    82901772.07797190546989441
    82901771.06932705640792847
     83217396.6076599508523941
    83217396.60766036808490753
    82901772.07797145843505859
    83217396.60766032338142395
    83217396.60766017436981201
    83217395.59517517685890198
    82901772.07797172665596008
    83217394.85398450493812561
     83217396.6076604425907135
    82901772.07797157764434814
    83217396.60765974223613739
    82901772.07797171175479889
    83217396.60765975713729858
    83217396.60766041278839111
    82901771.06932675838470459
    82901771.06932680308818817
    83217396.60766030848026276
    82901772.07797171175479889
    83217396.60766030848026276
    82901772.07797135412693024
     82901772.0779716819524765
    83217396.60766024887561798
    82901772.07797178626060486
    83217396.60766007006168365
    83217396.60765999555587769
    83217396.60765951871871948
    82901770.33094756305217743
    82901772.07797183096408844
    82901772.07797160744667053
    83217396.60766023397445679
    83217395.59517547488212585
    83217396.60765987634658813
     83217396.6076599657535553
    83217396.60766038298606873
    83217396.60765990614891052
    82901772.07797187566757202
    83217396.60766029357910156
    82901772.07797171175479889
    83217396.60766015946865082
    82901772.07797142863273621
    82901772.07797208428382874
    82901771.06932723522186279
    82901772.07797175645828247
    82901772.07797183096408844
    82901772.07797220349311829
    82901772.07797181606292725
    82901772.07797123491764069
    82901772.07797151803970337
    83217396.60766018927097321
     82901771.0693267434835434
    82901772.07797187566757202
    82901772.07797187566757202
    82901772.07797172665596008
    82901772.07797218859195709
     82901770.3309473842382431
    82901772.07797162234783173
    82901772.07797153294086456
    82901772.07797181606292725
    83217396.60766018927097321
    83217396.60766024887561798
    83217396.60765990614891052
    82901772.07797181606292725
    82901772.07797113060951233
    82901772.07797175645828247
    82901772.07797156274318695
    82901771.06932733952999115
    82901772.07797165215015411
    82901771.06932705640792847
    83217396.60766045749187469
     83217395.5951753556728363
    83217396.60766002535820007
     83217394.8539850264787674
    82901772.07797175645828247
    82901772.07797190546989441
    83217396.60766030848026276
    83217396.60765987634658813
!Field "H_inverse_eigen_max" Scalar 1
    83217396.60766057670116425
     82901772.0779714435338974
    82901772.07797203958034515
    83217396.60766021907329559
    83217398.63263022899627686
    83217396.60766038298606873
     82901772.0779716968536377
    83217398.36133569478988647
    82901772.07797181606292725
    83217396.60766029357910156
    82901774.09526163339614868
    83217396.60766001045703888
    82901773.82499583065509796
    82901772.07797202467918396
    82901772.07797145843505859
    83217396.60766048729419708
    83217398.63263051211833954
    83217396.60765953361988068
    82901772.07797208428382874
    83217396.60766023397445679
    83217396.60766036808490753
    83217396.60766047239303589
    82901772.07797190546989441
    82901774.09526176750659943
     83217396.6076599508523941
    83217396.60766036808490753
    82901772.07797145843505859
    83217396.60766032338142395
    83217396.60766017436981201
    83217398.63263025879859924
    82901772.07797172665596008
    83217398.36133551597595215
     83217396.6076604425907135
    82901772.07797157764434814
    83217396.60765974223613739
    82901772.07797171175479889
    83217396.60765975713729858
    83217396.60766041278839111
    82901774.09526145458221436
    82901774.09526151418685913
    83217396.60766030848026276
    82901772.07797171175479889
    83217396.60766030848026276
    82901772.07797135412693024
     82901772.0779716819524765
    83217396.60766024887561798
    82901772.07797178626060486
    83217396.60766007006168365
    83217396.60765999555587769
    83217396.60765951871871948
    82901773.82499599456787109
    82901772.07797183096408844
    82901772.07797160744667053
    83217396.60766023397445679
    83217398.63263055682182312
    83217396.60765987634658813
     83217396.6076599657535553
    83217396.60766038298606873
    83217396.60765990614891052
    82901772.07797187566757202
    83217396.60766029357910156
    82901772.07797171175479889
    83217396.60766015946865082
    82901772.07797142863273621
    82901772.07797208428382874
    82901774.09526194632053375
    82901772.07797175645828247
    82901772.07797183096408844
    82901772.07797220349311829
    82901772.07797181606292725
    82901772.07797123491764069
    82901772.07797151803970337
    83217396.60766018927097321
    82901774.09526145458221436
    82901772.07797187566757202
    82901772.07797187566757202
    82901772.07797172665596008
    82901772.07797218859195709
    82901773.82499581575393677
    82901772.07797162234783173
    82901772.07797153294086456
    82901772.07797181606292725
    83217396.60766018927097321
    83217396.60766024887561798
    83217396.60765990614891052
    82901772.07797181606292725
    82901772.07797113060951233
    82901772.07797175645828247
    82901772.07797156274318695
    82901774.09526203572750092
    82901772.07797165215015411
    82901774.09526176750659943
    83217396.60766045749187469
    83217398.63263042271137238
    83217396.60766002535820007
    83217398.36133603751659393
    82901772.07797175645828247
    82901772.07797190546989441
    83217396.60766030848026276
    83217396.60765987634658813
!Field "hmin" Scalar 1
    83217396.60766059160232544
    82901772.07797145843505859
    82901772.07797203958034515
    83217396.60766024887561798
    83217396.60766017436981201
    83217394.58269037306308746
    82901772.07797171175479889
    83217396.60766018927097321
    82901772.07797183096408844
     83217394.5826902836561203
    82901770.06068205833435059
    83217396.60766004025936127
    82901772.07797160744667053
    82901772.07797203958034515
    82901769.22509296238422394
    83217394.58269050717353821
    83217396.60766045749187469
    83217396.60765954852104187
    82901772.07797208428382874
    83217396.60766024887561798
    83217396.60766038298606873
    83217396.60766048729419708
     82901772.0779719203710556
    82901770.06068219244480133
     83217396.6076599508523941
    83217396.60766035318374634
    82901772.07797145843505859
    83217396.60766033828258514
    83217396.60766018927097321
    83217394.85398472845554352
    82901772.07797172665596008
    83217394.58268997073173523
    83217396.60766045749187469
    82901772.07797160744667053
    83217394.58268976211547852
    82901772.07797174155712128
    83217396.60765977203845978
    83217396.60766041278839111
    82901772.07797165215015411
    82901772.07797171175479889
    83217396.60766032338142395
    82901772.07797171175479889
    83217396.60766032338142395
    82901772.07797136902809143
    82901772.07797171175479889
    83217394.58269025385379791
    82901770.06068204343318939
    83217396.60766009986400604
    83217396.60765999555587769
    83217396.60765951871871948
    82901772.07797178626060486
    82901772.07797183096408844
    82901772.07797162234783173
    83217396.60766024887561798
    83217396.60766048729419708
    83217396.60765989124774933
     83217396.6076599657535553
    83217396.60766039788722992
    83217396.60765992105007172
    82901772.07797187566757202
    83217396.60766032338142395
    82901772.07797172665596008
    83217396.60766015946865082
    82901772.07797142863273621
    82901772.07797208428382874
     82901772.0779721587896347
    82901772.07797175645828247
    82901770.33094766736030579
    82901772.07797223329544067
    82901772.07797181606292725
    82901772.07797124981880188
    82901772.07797151803970337
     83217396.6076602041721344
    82901772.07797163724899292
    82901772.07797187566757202
    82901770.06068211793899536
    82901772.07797175645828247
    82901772.07797220349311829
    82901772.07797159254550934
    82901770.06068186461925507
    82901770.06068176031112671
    82901770.06068205833435059
    83217394.85398472845554352
    83217396.60766027867794037
    83217396.60765992105007172
    82901772.07797183096408844
    82901772.07797111570835114
    82901772.07797175645828247
    82901772.07797157764434814
    82901770.06068246066570282
    82901772.07797166705131531
    82901770.06068219244480133
     83217396.6076604425907135
    83217396.60766039788722992
    83217396.60766004025936127
    83217394.58269055187702179
    82901770.33094756305217743
    82901772.07797190546989441
    83217394.58269031345844269
    83217396.60765989124774933
!Field "hmax" Scalar 1
    83217396.60766059160232544
    82901772.07797145843505859
    82901772.07797203958034515
    83217396.60766024887561798
    83217396.60766017436981201
    83217397.62014542520046234
    82901772.07797171175479889
    83217396.60766018927097321
    82901772.07797183096408844
    83217397.62014532089233398
    82901773.08661672472953796
    83217396.60766004025936127
    82901772.07797160744667053
    82901772.07797203958034515
    82901773.50441078841686249
     83217397.6201455295085907
    83217396.60766045749187469
    83217396.60765954852104187
    82901772.07797208428382874
    83217396.60766024887561798
    83217396.60766038298606873
    83217396.60766048729419708
     82901772.0779719203710556
    82901773.08661685883998871
     83217396.6076599508523941
    83217396.60766035318374634
    82901772.07797145843505859
    83217396.60766033828258514
    83217396.60766018927097321
    83217398.36133575439453125
    82901772.07797172665596008
    83217397.62014502286911011
    83217396.60766045749187469
    82901772.07797160744667053
    83217397.62014478445053101
    82901772.07797174155712128
    83217396.60765977203845978
    83217396.60766041278839111
    82901772.07797165215015411
    82901772.07797171175479889
    83217396.60766032338142395
    82901772.07797171175479889
    83217396.60766032338142395
    82901772.07797136902809143
    82901772.07797171175479889
    83217397.62014530599117279
    82901773.08661670982837677
    83217396.60766009986400604
    83217396.60765999555587769
    83217396.60765951871871948
    82901772.07797178626060486
    82901772.07797183096408844
    82901772.07797162234783173
    83217396.60766024887561798
    83217396.60766048729419708
    83217396.60765989124774933
     83217396.6076599657535553
    83217396.60766039788722992
    83217396.60765992105007172
    82901772.07797187566757202
    83217396.60766032338142395
    82901772.07797172665596008
    83217396.60766015946865082
    82901772.07797142863273621
    82901772.07797208428382874
     82901772.0779721587896347
    82901772.07797175645828247
    82901773.82499608397483826
    82901772.07797223329544067
    82901772.07797181606292725
    82901772.07797124981880188
    82901772.07797151803970337
     83217396.6076602041721344
    82901772.07797163724899292
    82901772.07797187566757202
    82901773.08661678433418274
    82901772.07797175645828247
    82901772.07797220349311829
    82901772.07797159254550934
    82901773.08661653101444244
    82901773.08661644160747528
    82901773.08661672472953796
    83217398.36133575439453125
    83217396.60766027867794037
    83217396.60765992105007172
    82901772.07797183096408844
    82901772.07797111570835114
    82901772.07797175645828247
    82901772.07797157764434814
      82901773.086617112159729
    82901772.07797166705131531
    82901773.08661685883998871
     83217396.6076604425907135
    83217396.60766039788722992
    83217396.60766004025936127
    83217397.62014557421207428
    82901773.82499599456787109
    82901772.07797190546989441
    83217397.62014535069465637
    83217396.60765989124774933
!Field "hmin_hmax_ratio" Scalar 1
                             1
                             1
                             1
                             1
                             1
   0.9999999634997591702045838
                             1
                             1
                             1
   0.9999999634997592812268863
   0.9999999634997595032714912
                             1
                             1
                             1
    0.999999948380865144592633
   0.9999999634997593922491887
                             1
                             1
                             1
                             1
                             1
                             1
                             1
   0.9999999634997592812268863
                             1
                             1
                             1
                             1
                             1
   0.9999999578531523214408594
                             1
   0.9999999634997592812268863
                             1
                             1
   0.9999999634997593922491887
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
   0.9999999634997591702045838
   0.9999999634997592812268863
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
                             1
   0.9999999578531524324631619
                             1
                             1
                             1
                             1
                             1
                             1
                             1
   0.9999999634997592812268863
                             1
                             1
                             1
   0.9999999634997592812268863
   0.9999999634997592812268863
   0.9999999634997592812268863
   0.9999999578531523214408594
                             1
                             1
                             1
                             1
                             1
                             1
   0.9999999634997595032714912
                             1
   0.9999999634997595032714912
                             1
                             1
                             1
   0.9999999634997593922491887
   0.9999999578531524324631619
                             1
   0.9999999634997592812268863
                             1
!Field "Domains" Scalar 1
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
                             0
